magic
tech sky130A
magscale 1 2
timestamp 1654523691
<< viali >>
rect 10609 37349 10643 37383
rect 34161 37349 34195 37383
rect 9321 37281 9355 37315
rect 11989 37281 12023 37315
rect 14933 37281 14967 37315
rect 17233 37281 17267 37315
rect 20637 37281 20671 37315
rect 27261 37281 27295 37315
rect 32137 37281 32171 37315
rect 33517 37281 33551 37315
rect 36737 37281 36771 37315
rect 1409 37213 1443 37247
rect 2329 37213 2363 37247
rect 2973 37213 3007 37247
rect 5641 37213 5675 37247
rect 6653 37213 6687 37247
rect 7297 37213 7331 37247
rect 7757 37213 7791 37247
rect 9781 37213 9815 37247
rect 11529 37213 11563 37247
rect 14105 37213 14139 37247
rect 17693 37213 17727 37247
rect 18705 37213 18739 37247
rect 19441 37213 19475 37247
rect 21833 37213 21867 37247
rect 23029 37213 23063 37247
rect 23673 37213 23707 37247
rect 24409 37213 24443 37247
rect 25421 37213 25455 37247
rect 25881 37213 25915 37247
rect 26985 37213 27019 37247
rect 29745 37213 29779 37247
rect 34897 37213 34931 37247
rect 37289 37213 37323 37247
rect 37933 37213 37967 37247
rect 3801 37145 3835 37179
rect 5457 37145 5491 37179
rect 7205 37145 7239 37179
rect 11713 37145 11747 37179
rect 19625 37145 19659 37179
rect 29929 37145 29963 37179
rect 31585 37145 31619 37179
rect 35081 37145 35115 37179
rect 38025 37145 38059 37179
rect 1593 37077 1627 37111
rect 2237 37077 2271 37111
rect 2881 37077 2915 37111
rect 6469 37077 6503 37111
rect 14197 37077 14231 37111
rect 21925 37077 21959 37111
rect 22937 37077 22971 37111
rect 25973 37077 26007 37111
rect 28733 37077 28767 37111
rect 37381 37077 37415 37111
rect 10885 36873 10919 36907
rect 1593 36805 1627 36839
rect 3249 36805 3283 36839
rect 3893 36805 3927 36839
rect 14289 36805 14323 36839
rect 21833 36805 21867 36839
rect 28549 36805 28583 36839
rect 29285 36805 29319 36839
rect 35081 36805 35115 36839
rect 37473 36805 37507 36839
rect 5733 36737 5767 36771
rect 6469 36737 6503 36771
rect 7205 36737 7239 36771
rect 10793 36737 10827 36771
rect 11529 36737 11563 36771
rect 16129 36737 16163 36771
rect 17141 36737 17175 36771
rect 17693 36737 17727 36771
rect 21189 36737 21223 36771
rect 23673 36737 23707 36771
rect 24133 36737 24167 36771
rect 27813 36737 27847 36771
rect 28457 36737 28491 36771
rect 34897 36737 34931 36771
rect 36737 36737 36771 36771
rect 37381 36737 37415 36771
rect 3433 36669 3467 36703
rect 5549 36669 5583 36703
rect 8401 36669 8435 36703
rect 8585 36669 8619 36703
rect 9781 36669 9815 36703
rect 11713 36669 11747 36703
rect 11989 36669 12023 36703
rect 15945 36669 15979 36703
rect 17877 36669 17911 36703
rect 18153 36669 18187 36703
rect 20729 36669 20763 36703
rect 23489 36669 23523 36703
rect 24317 36669 24351 36703
rect 24593 36669 24627 36703
rect 29101 36669 29135 36703
rect 30481 36669 30515 36703
rect 32413 36669 32447 36703
rect 32597 36669 32631 36703
rect 32873 36669 32907 36703
rect 17049 36533 17083 36567
rect 27353 36533 27387 36567
rect 27905 36533 27939 36567
rect 31585 36533 31619 36567
rect 9045 36329 9079 36363
rect 17049 36329 17083 36363
rect 17877 36329 17911 36363
rect 24501 36329 24535 36363
rect 29653 36329 29687 36363
rect 30205 36329 30239 36363
rect 34805 36329 34839 36363
rect 1409 36193 1443 36227
rect 3065 36193 3099 36227
rect 4629 36193 4663 36227
rect 5825 36193 5859 36227
rect 7757 36193 7791 36227
rect 9781 36193 9815 36227
rect 10333 36193 10367 36227
rect 19257 36193 19291 36227
rect 19993 36193 20027 36227
rect 25789 36193 25823 36227
rect 25973 36193 26007 36227
rect 26433 36193 26467 36227
rect 31677 36193 31711 36227
rect 32229 36193 32263 36227
rect 38117 36193 38151 36227
rect 3249 36125 3283 36159
rect 6469 36125 6503 36159
rect 9137 36125 9171 36159
rect 12173 36125 12207 36159
rect 13001 36125 13035 36159
rect 15853 36125 15887 36159
rect 16497 36125 16531 36159
rect 17141 36125 17175 36159
rect 17785 36125 17819 36159
rect 18521 36125 18555 36159
rect 21557 36125 21591 36159
rect 23029 36125 23063 36159
rect 24593 36125 24627 36159
rect 25237 36125 25271 36159
rect 28457 36125 28491 36159
rect 28641 36125 28675 36159
rect 29561 36125 29595 36159
rect 34161 36125 34195 36159
rect 34713 36125 34747 36159
rect 35817 36125 35851 36159
rect 36277 36125 36311 36159
rect 5641 36057 5675 36091
rect 7113 36057 7147 36091
rect 9965 36057 9999 36091
rect 12265 36057 12299 36091
rect 13185 36057 13219 36091
rect 15577 36057 15611 36091
rect 18613 36057 18647 36091
rect 19441 36057 19475 36091
rect 22385 36057 22419 36091
rect 31861 36057 31895 36091
rect 36461 36057 36495 36091
rect 12817 35989 12851 36023
rect 14105 35989 14139 36023
rect 16313 35989 16347 36023
rect 25145 35989 25179 36023
rect 28549 35989 28583 36023
rect 4537 35785 4571 35819
rect 9781 35785 9815 35819
rect 10425 35785 10459 35819
rect 14841 35785 14875 35819
rect 21925 35785 21959 35819
rect 27169 35785 27203 35819
rect 30205 35785 30239 35819
rect 32229 35785 32263 35819
rect 32873 35785 32907 35819
rect 37473 35785 37507 35819
rect 5365 35717 5399 35751
rect 14565 35717 14599 35751
rect 16037 35717 16071 35751
rect 35081 35717 35115 35751
rect 36737 35717 36771 35751
rect 4629 35649 4663 35683
rect 5733 35649 5767 35683
rect 6469 35649 6503 35683
rect 8401 35649 8435 35683
rect 9689 35649 9723 35683
rect 10517 35649 10551 35683
rect 14197 35649 14231 35683
rect 14355 35649 14389 35683
rect 14473 35649 14507 35683
rect 14657 35649 14691 35683
rect 15301 35649 15335 35683
rect 15485 35649 15519 35683
rect 15945 35649 15979 35683
rect 17049 35649 17083 35683
rect 19533 35649 19567 35683
rect 20453 35649 20487 35683
rect 22017 35649 22051 35683
rect 22661 35649 22695 35683
rect 25329 35649 25363 35683
rect 26157 35649 26191 35683
rect 27353 35649 27387 35683
rect 27813 35649 27847 35683
rect 30113 35649 30147 35683
rect 32321 35649 32355 35683
rect 32965 35649 32999 35683
rect 34897 35649 34931 35683
rect 37381 35649 37415 35683
rect 1777 35581 1811 35615
rect 1961 35581 1995 35615
rect 2789 35581 2823 35615
rect 7205 35581 7239 35615
rect 11713 35581 11747 35615
rect 11989 35581 12023 35615
rect 17325 35581 17359 35615
rect 20821 35581 20855 35615
rect 22845 35581 22879 35615
rect 23213 35581 23247 35615
rect 27997 35581 28031 35615
rect 28365 35581 28399 35615
rect 15301 35513 15335 35547
rect 19717 35513 19751 35547
rect 13461 35445 13495 35479
rect 18797 35445 18831 35479
rect 25145 35445 25179 35479
rect 26065 35445 26099 35479
rect 4077 35241 4111 35275
rect 12265 35241 12299 35275
rect 13461 35241 13495 35275
rect 17693 35241 17727 35275
rect 19349 35241 19383 35275
rect 27353 35241 27387 35275
rect 29561 35241 29595 35275
rect 32413 35241 32447 35275
rect 28825 35173 28859 35207
rect 2697 35105 2731 35139
rect 12909 35105 12943 35139
rect 15117 35105 15151 35139
rect 15669 35105 15703 35139
rect 17049 35105 17083 35139
rect 24869 35105 24903 35139
rect 27721 35105 27755 35139
rect 31033 35105 31067 35139
rect 37197 35105 37231 35139
rect 3249 35037 3283 35071
rect 3985 35037 4019 35071
rect 5825 35037 5859 35071
rect 6469 35037 6503 35071
rect 8953 35037 8987 35071
rect 11253 35037 11287 35071
rect 11529 35037 11563 35071
rect 12449 35037 12483 35071
rect 13369 35037 13403 35071
rect 13553 35037 13587 35071
rect 14289 35037 14323 35071
rect 15485 35037 15519 35071
rect 16405 35037 16439 35071
rect 16589 35037 16623 35071
rect 17509 35037 17543 35071
rect 18521 35037 18555 35071
rect 19441 35037 19475 35071
rect 20729 35037 20763 35071
rect 23857 35037 23891 35071
rect 27537 35037 27571 35071
rect 28273 35037 28307 35071
rect 28549 35037 28583 35071
rect 28641 35037 28675 35071
rect 31309 35037 31343 35071
rect 35817 35037 35851 35071
rect 38117 35037 38151 35071
rect 3065 34969 3099 35003
rect 5457 34969 5491 35003
rect 6837 34969 6871 35003
rect 9229 34969 9263 35003
rect 11345 34969 11379 35003
rect 12541 34969 12575 35003
rect 12633 34969 12667 35003
rect 12771 34969 12805 35003
rect 15393 34969 15427 35003
rect 17187 34969 17221 35003
rect 17325 34969 17359 35003
rect 17417 34969 17451 35003
rect 18153 34969 18187 35003
rect 18337 34969 18371 35003
rect 21373 34969 21407 35003
rect 25145 34969 25179 35003
rect 28457 34969 28491 35003
rect 37933 34969 37967 35003
rect 10701 34901 10735 34935
rect 11713 34901 11747 34935
rect 14197 34901 14231 34935
rect 15301 34901 15335 34935
rect 16589 34901 16623 34935
rect 23673 34901 23707 34935
rect 26617 34901 26651 34935
rect 2237 34697 2271 34731
rect 2881 34697 2915 34731
rect 10793 34697 10827 34731
rect 13001 34697 13035 34731
rect 15117 34697 15151 34731
rect 17141 34697 17175 34731
rect 17969 34697 18003 34731
rect 22293 34697 22327 34731
rect 25513 34697 25547 34731
rect 27997 34697 28031 34731
rect 29009 34697 29043 34731
rect 37565 34697 37599 34731
rect 11529 34629 11563 34663
rect 11897 34629 11931 34663
rect 12035 34629 12069 34663
rect 12633 34629 12667 34663
rect 12849 34629 12883 34663
rect 14473 34629 14507 34663
rect 23581 34629 23615 34663
rect 27169 34629 27203 34663
rect 27385 34629 27419 34663
rect 28549 34629 28583 34663
rect 32229 34629 32263 34663
rect 36553 34629 36587 34663
rect 1685 34561 1719 34595
rect 2329 34561 2363 34595
rect 2973 34561 3007 34595
rect 10885 34561 10919 34595
rect 11713 34561 11747 34595
rect 11805 34561 11839 34595
rect 12173 34561 12207 34595
rect 14013 34561 14047 34595
rect 15394 34561 15428 34595
rect 15577 34561 15611 34595
rect 17233 34561 17267 34595
rect 17785 34561 17819 34595
rect 18981 34561 19015 34595
rect 20085 34561 20119 34595
rect 21189 34561 21223 34595
rect 22477 34561 22511 34595
rect 23305 34561 23339 34595
rect 25881 34561 25915 34595
rect 28181 34561 28215 34595
rect 28273 34561 28307 34595
rect 28365 34561 28399 34595
rect 29285 34561 29319 34595
rect 29837 34561 29871 34595
rect 32321 34561 32355 34595
rect 33425 34561 33459 34595
rect 36737 34561 36771 34595
rect 37473 34561 37507 34595
rect 3617 34493 3651 34527
rect 3801 34493 3835 34527
rect 4169 34493 4203 34527
rect 8493 34493 8527 34527
rect 14197 34493 14231 34527
rect 15301 34493 15335 34527
rect 15485 34493 15519 34527
rect 20913 34493 20947 34527
rect 25053 34493 25087 34527
rect 25973 34493 26007 34527
rect 26157 34493 26191 34527
rect 29009 34493 29043 34527
rect 33793 34493 33827 34527
rect 35817 34493 35851 34527
rect 27537 34425 27571 34459
rect 29193 34425 29227 34459
rect 8756 34357 8790 34391
rect 10241 34357 10275 34391
rect 12817 34357 12851 34391
rect 13829 34357 13863 34391
rect 14381 34357 14415 34391
rect 18889 34357 18923 34391
rect 19993 34357 20027 34391
rect 27353 34357 27387 34391
rect 30100 34357 30134 34391
rect 31585 34357 31619 34391
rect 1961 34153 1995 34187
rect 3893 34153 3927 34187
rect 9873 34153 9907 34187
rect 11713 34153 11747 34187
rect 14289 34153 14323 34187
rect 17141 34153 17175 34187
rect 25237 34153 25271 34187
rect 29929 34153 29963 34187
rect 2605 34085 2639 34119
rect 18429 34085 18463 34119
rect 3249 34017 3283 34051
rect 10977 34017 11011 34051
rect 11253 34017 11287 34051
rect 15393 34017 15427 34051
rect 18337 34017 18371 34051
rect 18705 34017 18739 34051
rect 20729 34017 20763 34051
rect 21925 34017 21959 34051
rect 25605 34017 25639 34051
rect 27905 34017 27939 34051
rect 27997 34017 28031 34051
rect 37381 34017 37415 34051
rect 3985 33949 4019 33983
rect 4445 33949 4479 33983
rect 5365 33949 5399 33983
rect 6653 33949 6687 33983
rect 9965 33949 9999 33983
rect 10885 33949 10919 33983
rect 11897 33949 11931 33983
rect 11989 33949 12023 33983
rect 12265 33949 12299 33983
rect 13001 33949 13035 33983
rect 13093 33949 13127 33983
rect 13277 33949 13311 33983
rect 13369 33949 13403 33983
rect 18245 33949 18279 33983
rect 18521 33949 18555 33983
rect 21005 33949 21039 33983
rect 21649 33949 21683 33983
rect 24593 33949 24627 33983
rect 24685 33949 24719 33983
rect 25421 33949 25455 33983
rect 26065 33949 26099 33983
rect 26249 33949 26283 33983
rect 26433 33949 26467 33983
rect 27077 33949 27111 33983
rect 27721 33949 27755 33983
rect 27813 33949 27847 33983
rect 29837 33949 29871 33983
rect 30665 33949 30699 33983
rect 32045 33949 32079 33983
rect 36277 33949 36311 33983
rect 6009 33881 6043 33915
rect 7481 33881 7515 33915
rect 12081 33881 12115 33915
rect 14257 33881 14291 33915
rect 14473 33881 14507 33915
rect 15669 33881 15703 33915
rect 32321 33881 32355 33915
rect 36461 33881 36495 33915
rect 4629 33813 4663 33847
rect 12817 33813 12851 33847
rect 14105 33813 14139 33847
rect 19257 33813 19291 33847
rect 23397 33813 23431 33847
rect 24409 33813 24443 33847
rect 26893 33813 26927 33847
rect 27537 33813 27571 33847
rect 30573 33813 30607 33847
rect 33793 33813 33827 33847
rect 15761 33609 15795 33643
rect 16957 33609 16991 33643
rect 18521 33609 18555 33643
rect 22937 33609 22971 33643
rect 23305 33609 23339 33643
rect 24961 33609 24995 33643
rect 25789 33609 25823 33643
rect 27629 33609 27663 33643
rect 33241 33609 33275 33643
rect 37381 33609 37415 33643
rect 9781 33541 9815 33575
rect 11713 33541 11747 33575
rect 15393 33541 15427 33575
rect 17969 33541 18003 33575
rect 22201 33541 22235 33575
rect 23397 33541 23431 33575
rect 30481 33541 30515 33575
rect 2145 33473 2179 33507
rect 3617 33473 3651 33507
rect 4997 33473 5031 33507
rect 8401 33473 8435 33507
rect 9045 33473 9079 33507
rect 9873 33473 9907 33507
rect 10333 33473 10367 33507
rect 10609 33473 10643 33507
rect 17049 33473 17083 33507
rect 18061 33473 18095 33507
rect 18889 33473 18923 33507
rect 21281 33473 21315 33507
rect 22477 33473 22511 33507
rect 24501 33473 24535 33507
rect 25605 33473 25639 33507
rect 26985 33473 27019 33507
rect 27905 33473 27939 33507
rect 28089 33473 28123 33507
rect 32137 33473 32171 33507
rect 33333 33473 33367 33507
rect 36553 33473 36587 33507
rect 37473 33473 37507 33507
rect 38117 33473 38151 33507
rect 5365 33405 5399 33439
rect 10425 33405 10459 33439
rect 12633 33405 12667 33439
rect 12909 33405 12943 33439
rect 14381 33405 14415 33439
rect 15117 33405 15151 33439
rect 15301 33405 15335 33439
rect 17601 33405 17635 33439
rect 18705 33405 18739 33439
rect 18797 33405 18831 33439
rect 18981 33405 19015 33439
rect 19533 33405 19567 33439
rect 21005 33405 21039 33439
rect 22201 33405 22235 33439
rect 23489 33405 23523 33439
rect 24593 33405 24627 33439
rect 24685 33405 24719 33439
rect 24780 33405 24814 33439
rect 25421 33405 25455 33439
rect 27813 33405 27847 33439
rect 27997 33405 28031 33439
rect 30757 33405 30791 33439
rect 11529 33337 11563 33371
rect 8493 33269 8527 33303
rect 9137 33269 9171 33303
rect 10333 33269 10367 33303
rect 10793 33269 10827 33303
rect 17785 33269 17819 33303
rect 22385 33269 22419 33303
rect 27077 33269 27111 33303
rect 29009 33269 29043 33303
rect 32321 33269 32355 33303
rect 8953 33065 8987 33099
rect 12817 33065 12851 33099
rect 14841 33065 14875 33099
rect 18429 33065 18463 33099
rect 20729 33065 20763 33099
rect 22753 33065 22787 33099
rect 23581 33065 23615 33099
rect 24685 33065 24719 33099
rect 27813 33065 27847 33099
rect 28641 33065 28675 33099
rect 30205 33065 30239 33099
rect 30665 33065 30699 33099
rect 31769 33065 31803 33099
rect 19809 32997 19843 33031
rect 7573 32929 7607 32963
rect 10701 32929 10735 32963
rect 13001 32929 13035 32963
rect 13461 32929 13495 32963
rect 15485 32929 15519 32963
rect 18337 32929 18371 32963
rect 26065 32929 26099 32963
rect 26341 32929 26375 32963
rect 31953 32929 31987 32963
rect 32137 32929 32171 32963
rect 5825 32861 5859 32895
rect 7757 32861 7791 32895
rect 7849 32861 7883 32895
rect 11345 32861 11379 32895
rect 11437 32861 11471 32895
rect 11621 32861 11655 32895
rect 11713 32861 11747 32895
rect 12173 32861 12207 32895
rect 13093 32861 13127 32895
rect 14289 32861 14323 32895
rect 14933 32861 14967 32895
rect 18521 32861 18555 32895
rect 19257 32861 19291 32895
rect 19533 32861 19567 32895
rect 19625 32861 19659 32895
rect 20821 32861 20855 32895
rect 21373 32861 21407 32895
rect 22661 32861 22695 32895
rect 25421 32861 25455 32895
rect 28641 32861 28675 32895
rect 28733 32861 28767 32895
rect 29929 32861 29963 32895
rect 30021 32861 30055 32895
rect 30849 32861 30883 32895
rect 31033 32861 31067 32895
rect 31171 32861 31205 32895
rect 31309 32861 31343 32895
rect 32045 32861 32079 32895
rect 32229 32861 32263 32895
rect 32781 32861 32815 32895
rect 33977 32861 34011 32895
rect 34713 32861 34747 32895
rect 36277 32861 36311 32895
rect 5273 32793 5307 32827
rect 10425 32793 10459 32827
rect 12265 32793 12299 32827
rect 13369 32793 13403 32827
rect 15761 32793 15795 32827
rect 18245 32793 18279 32827
rect 19441 32793 19475 32827
rect 21741 32793 21775 32827
rect 23765 32793 23799 32827
rect 24869 32793 24903 32827
rect 30941 32793 30975 32827
rect 32965 32793 32999 32827
rect 33793 32793 33827 32827
rect 36461 32793 36495 32827
rect 38117 32793 38151 32827
rect 7573 32725 7607 32759
rect 11161 32725 11195 32759
rect 14197 32725 14231 32759
rect 17233 32725 17267 32759
rect 18705 32725 18739 32759
rect 23397 32725 23431 32759
rect 23565 32725 23599 32759
rect 24501 32725 24535 32759
rect 24669 32725 24703 32759
rect 25513 32725 25547 32759
rect 29009 32725 29043 32759
rect 29561 32725 29595 32759
rect 33149 32725 33183 32759
rect 34161 32725 34195 32759
rect 34805 32725 34839 32759
rect 11529 32521 11563 32555
rect 13093 32521 13127 32555
rect 15209 32521 15243 32555
rect 17969 32521 18003 32555
rect 21281 32521 21315 32555
rect 25329 32521 25363 32555
rect 26249 32521 26283 32555
rect 27797 32521 27831 32555
rect 28625 32521 28659 32555
rect 30113 32521 30147 32555
rect 31033 32521 31067 32555
rect 31217 32521 31251 32555
rect 32229 32521 32263 32555
rect 35173 32521 35207 32555
rect 37657 32521 37691 32555
rect 10241 32453 10275 32487
rect 11897 32453 11931 32487
rect 13185 32453 13219 32487
rect 13829 32453 13863 32487
rect 14565 32453 14599 32487
rect 15485 32453 15519 32487
rect 19073 32453 19107 32487
rect 22109 32453 22143 32487
rect 27997 32453 28031 32487
rect 28825 32453 28859 32487
rect 29745 32453 29779 32487
rect 30849 32453 30883 32487
rect 31125 32453 31159 32487
rect 32505 32453 32539 32487
rect 5825 32385 5859 32419
rect 6837 32385 6871 32419
rect 7021 32385 7055 32419
rect 9965 32385 9999 32419
rect 10793 32385 10827 32419
rect 11713 32385 11747 32419
rect 11805 32385 11839 32419
rect 12035 32385 12069 32419
rect 14013 32385 14047 32419
rect 15393 32385 15427 32419
rect 15577 32385 15611 32419
rect 15761 32385 15795 32419
rect 17049 32385 17083 32419
rect 17877 32385 17911 32419
rect 18889 32385 18923 32419
rect 19257 32385 19291 32419
rect 19717 32385 19751 32419
rect 21097 32385 21131 32419
rect 21833 32385 21867 32419
rect 24409 32385 24443 32419
rect 25605 32385 25639 32419
rect 26065 32385 26099 32419
rect 26985 32385 27019 32419
rect 27169 32385 27203 32419
rect 29653 32385 29687 32419
rect 29929 32385 29963 32419
rect 31401 32385 31435 32419
rect 32413 32385 32447 32419
rect 32597 32385 32631 32419
rect 32735 32385 32769 32419
rect 36553 32385 36587 32419
rect 37749 32385 37783 32419
rect 7481 32317 7515 32351
rect 7757 32317 7791 32351
rect 9873 32317 9907 32351
rect 10333 32317 10367 32351
rect 12173 32317 12207 32351
rect 16957 32317 16991 32351
rect 19809 32317 19843 32351
rect 23581 32317 23615 32351
rect 24225 32317 24259 32351
rect 24317 32317 24351 32351
rect 24501 32317 24535 32351
rect 25329 32317 25363 32351
rect 32873 32317 32907 32351
rect 33425 32317 33459 32351
rect 33701 32317 33735 32351
rect 9689 32249 9723 32283
rect 16681 32249 16715 32283
rect 25513 32249 25547 32283
rect 27629 32249 27663 32283
rect 28457 32249 28491 32283
rect 1961 32181 1995 32215
rect 5733 32181 5767 32215
rect 6837 32181 6871 32215
rect 9229 32181 9263 32215
rect 10977 32181 11011 32215
rect 14657 32181 14691 32215
rect 24041 32181 24075 32215
rect 26985 32181 27019 32215
rect 27813 32181 27847 32215
rect 28641 32181 28675 32215
rect 36093 32181 36127 32215
rect 10609 31977 10643 32011
rect 12449 31977 12483 32011
rect 13277 31977 13311 32011
rect 18521 31977 18555 32011
rect 21005 31977 21039 32011
rect 22569 31977 22603 32011
rect 31401 31977 31435 32011
rect 7113 31909 7147 31943
rect 8401 31909 8435 31943
rect 14197 31909 14231 31943
rect 17233 31909 17267 31943
rect 24961 31909 24995 31943
rect 32229 31909 32263 31943
rect 1409 31841 1443 31875
rect 3249 31841 3283 31875
rect 6285 31841 6319 31875
rect 7297 31841 7331 31875
rect 8953 31841 8987 31875
rect 9321 31841 9355 31875
rect 11345 31841 11379 31875
rect 15577 31841 15611 31875
rect 17785 31841 17819 31875
rect 19257 31841 19291 31875
rect 22017 31841 22051 31875
rect 23029 31841 23063 31875
rect 23213 31841 23247 31875
rect 28733 31841 28767 31875
rect 29009 31841 29043 31875
rect 30481 31841 30515 31875
rect 32597 31841 32631 31875
rect 33517 31841 33551 31875
rect 34161 31841 34195 31875
rect 34713 31841 34747 31875
rect 34989 31841 35023 31875
rect 36277 31841 36311 31875
rect 6561 31773 6595 31807
rect 7389 31773 7423 31807
rect 7665 31773 7699 31807
rect 7757 31773 7791 31807
rect 8217 31773 8251 31807
rect 9137 31773 9171 31807
rect 10241 31773 10275 31807
rect 11069 31773 11103 31807
rect 12357 31773 12391 31807
rect 12541 31773 12575 31807
rect 13461 31773 13495 31807
rect 14105 31773 14139 31807
rect 14289 31773 14323 31807
rect 15301 31773 15335 31807
rect 16313 31773 16347 31807
rect 16497 31773 16531 31807
rect 17049 31773 17083 31807
rect 17693 31773 17727 31807
rect 17877 31773 17911 31807
rect 21925 31773 21959 31807
rect 22109 31773 22143 31807
rect 24685 31773 24719 31807
rect 25421 31773 25455 31807
rect 26157 31773 26191 31807
rect 27353 31773 27387 31807
rect 27721 31773 27755 31807
rect 29745 31773 29779 31807
rect 30573 31773 30607 31807
rect 31033 31773 31067 31807
rect 31401 31773 31435 31807
rect 31677 31773 31711 31807
rect 32413 31773 32447 31807
rect 33655 31773 33689 31807
rect 33977 31773 34011 31807
rect 38117 31773 38151 31807
rect 3065 31705 3099 31739
rect 10425 31705 10459 31739
rect 18505 31705 18539 31739
rect 18705 31705 18739 31739
rect 19533 31705 19567 31739
rect 22937 31705 22971 31739
rect 24409 31705 24443 31739
rect 24593 31705 24627 31739
rect 24777 31705 24811 31739
rect 27537 31705 27571 31739
rect 33793 31705 33827 31739
rect 33885 31705 33919 31739
rect 36461 31705 36495 31739
rect 4813 31637 4847 31671
rect 18337 31637 18371 31671
rect 25605 31637 25639 31671
rect 26341 31637 26375 31671
rect 29837 31637 29871 31671
rect 31217 31637 31251 31671
rect 2145 31433 2179 31467
rect 5733 31433 5767 31467
rect 10241 31433 10275 31467
rect 10409 31433 10443 31467
rect 17693 31433 17727 31467
rect 19257 31433 19291 31467
rect 20637 31433 20671 31467
rect 22293 31433 22327 31467
rect 23305 31433 23339 31467
rect 24225 31433 24259 31467
rect 24409 31433 24443 31467
rect 25237 31433 25271 31467
rect 32137 31433 32171 31467
rect 32965 31433 32999 31467
rect 33885 31433 33919 31467
rect 36645 31433 36679 31467
rect 7665 31365 7699 31399
rect 9413 31365 9447 31399
rect 9613 31365 9647 31399
rect 10609 31365 10643 31399
rect 11529 31365 11563 31399
rect 11729 31365 11763 31399
rect 14749 31365 14783 31399
rect 19809 31365 19843 31399
rect 24593 31365 24627 31399
rect 26985 31365 27019 31399
rect 32229 31365 32263 31399
rect 2237 31297 2271 31331
rect 5181 31297 5215 31331
rect 5641 31297 5675 31331
rect 5825 31297 5859 31331
rect 6653 31297 6687 31331
rect 7757 31297 7791 31331
rect 7849 31297 7883 31331
rect 8953 31297 8987 31331
rect 12357 31297 12391 31331
rect 15485 31297 15519 31331
rect 15669 31297 15703 31331
rect 17141 31297 17175 31331
rect 17877 31297 17911 31331
rect 18061 31297 18095 31331
rect 18153 31297 18187 31331
rect 18613 31297 18647 31331
rect 18981 31297 19015 31331
rect 19073 31297 19107 31331
rect 19901 31297 19935 31331
rect 20729 31297 20763 31331
rect 22385 31297 22419 31331
rect 23213 31297 23247 31331
rect 24041 31297 24075 31331
rect 24317 31297 24351 31331
rect 25053 31297 25087 31331
rect 26341 31297 26375 31331
rect 27169 31297 27203 31331
rect 27997 31297 28031 31331
rect 28365 31297 28399 31331
rect 31401 31297 31435 31331
rect 31585 31297 31619 31331
rect 32137 31297 32171 31331
rect 32413 31297 32447 31331
rect 33057 31297 33091 31331
rect 33793 31297 33827 31331
rect 33977 31297 34011 31331
rect 34621 31297 34655 31331
rect 36737 31297 36771 31331
rect 37657 31297 37691 31331
rect 12633 31229 12667 31263
rect 18705 31229 18739 31263
rect 23489 31229 23523 31263
rect 27905 31229 27939 31263
rect 30665 31229 30699 31263
rect 30941 31229 30975 31263
rect 6837 31161 6871 31195
rect 7481 31161 7515 31195
rect 8769 31161 8803 31195
rect 9781 31161 9815 31195
rect 14565 31161 14599 31195
rect 16957 31161 16991 31195
rect 26157 31161 26191 31195
rect 5089 31093 5123 31127
rect 8033 31093 8067 31127
rect 9597 31093 9631 31127
rect 10425 31093 10459 31127
rect 11713 31093 11747 31127
rect 11897 31093 11931 31127
rect 14105 31093 14139 31127
rect 15301 31093 15335 31127
rect 22845 31093 22879 31127
rect 27353 31093 27387 31127
rect 28365 31093 28399 31127
rect 28549 31093 28583 31127
rect 29193 31093 29227 31127
rect 31585 31093 31619 31127
rect 34529 31093 34563 31127
rect 35449 31093 35483 31127
rect 36093 31093 36127 31127
rect 37565 31093 37599 31127
rect 8217 30889 8251 30923
rect 9505 30889 9539 30923
rect 9689 30889 9723 30923
rect 10609 30889 10643 30923
rect 11069 30889 11103 30923
rect 23673 30889 23707 30923
rect 29561 30889 29595 30923
rect 7573 30821 7607 30855
rect 16221 30821 16255 30855
rect 17601 30821 17635 30855
rect 6101 30753 6135 30787
rect 10793 30753 10827 30787
rect 11529 30753 11563 30787
rect 12633 30753 12667 30787
rect 18153 30753 18187 30787
rect 18613 30753 18647 30787
rect 21465 30753 21499 30787
rect 27169 30753 27203 30787
rect 28641 30753 28675 30787
rect 36277 30753 36311 30787
rect 36461 30753 36495 30787
rect 7205 30685 7239 30719
rect 10885 30685 10919 30719
rect 11713 30685 11747 30719
rect 12817 30685 12851 30719
rect 12909 30685 12943 30719
rect 13001 30685 13035 30719
rect 13277 30685 13311 30719
rect 14473 30685 14507 30719
rect 16865 30685 16899 30719
rect 17417 30685 17451 30719
rect 18245 30685 18279 30719
rect 19717 30685 19751 30719
rect 21925 30685 21959 30719
rect 24777 30685 24811 30719
rect 28457 30685 28491 30719
rect 29745 30685 29779 30719
rect 29929 30685 29963 30719
rect 30113 30685 30147 30719
rect 31309 30685 31343 30719
rect 33793 30685 33827 30719
rect 35265 30685 35299 30719
rect 5825 30617 5859 30651
rect 7021 30617 7055 30651
rect 7297 30617 7331 30651
rect 8185 30617 8219 30651
rect 8401 30617 8435 30651
rect 9873 30617 9907 30651
rect 10609 30617 10643 30651
rect 13119 30617 13153 30651
rect 14749 30617 14783 30651
rect 19993 30617 20027 30651
rect 22201 30617 22235 30651
rect 26893 30617 26927 30651
rect 28365 30617 28399 30651
rect 29837 30617 29871 30651
rect 30573 30617 30607 30651
rect 30757 30617 30791 30651
rect 31493 30617 31527 30651
rect 33517 30617 33551 30651
rect 38117 30617 38151 30651
rect 4353 30549 4387 30583
rect 7389 30549 7423 30583
rect 8033 30549 8067 30583
rect 9673 30549 9707 30583
rect 11897 30549 11931 30583
rect 16681 30549 16715 30583
rect 24869 30549 24903 30583
rect 25421 30549 25455 30583
rect 28089 30549 28123 30583
rect 28273 30549 28307 30583
rect 32045 30549 32079 30583
rect 35357 30549 35391 30583
rect 7849 30345 7883 30379
rect 10425 30345 10459 30379
rect 12817 30345 12851 30379
rect 14289 30345 14323 30379
rect 14933 30345 14967 30379
rect 19717 30345 19751 30379
rect 22385 30345 22419 30379
rect 5365 30277 5399 30311
rect 8125 30277 8159 30311
rect 13277 30277 13311 30311
rect 13493 30277 13527 30311
rect 15209 30277 15243 30311
rect 15419 30277 15453 30311
rect 17049 30277 17083 30311
rect 20913 30277 20947 30311
rect 23121 30277 23155 30311
rect 25973 30277 26007 30311
rect 26985 30277 27019 30311
rect 27261 30277 27295 30311
rect 27471 30277 27505 30311
rect 28181 30277 28215 30311
rect 29009 30277 29043 30311
rect 33793 30277 33827 30311
rect 34529 30277 34563 30311
rect 4905 30209 4939 30243
rect 5641 30209 5675 30243
rect 6837 30209 6871 30243
rect 8033 30209 8067 30243
rect 8217 30209 8251 30243
rect 8401 30209 8435 30243
rect 9965 30209 9999 30243
rect 10241 30209 10275 30243
rect 11529 30209 11563 30243
rect 11621 30209 11655 30243
rect 12357 30209 12391 30243
rect 12632 30209 12666 30243
rect 14197 30209 14231 30243
rect 14473 30209 14507 30243
rect 15117 30209 15151 30243
rect 15301 30209 15335 30243
rect 16957 30209 16991 30243
rect 17141 30209 17175 30243
rect 18429 30209 18463 30243
rect 18705 30209 18739 30243
rect 19165 30209 19199 30243
rect 19349 30209 19383 30243
rect 19441 30209 19475 30243
rect 19533 30209 19567 30243
rect 20177 30209 20211 30243
rect 21005 30209 21039 30243
rect 22569 30209 22603 30243
rect 23213 30209 23247 30243
rect 23857 30209 23891 30243
rect 27170 30231 27204 30265
rect 27353 30209 27387 30243
rect 28089 30209 28123 30243
rect 28917 30209 28951 30243
rect 29101 30209 29135 30243
rect 29837 30209 29871 30243
rect 32229 30209 32263 30243
rect 33609 30209 33643 30243
rect 36461 30209 36495 30243
rect 37565 30209 37599 30243
rect 5549 30141 5583 30175
rect 6561 30141 6595 30175
rect 10057 30141 10091 30175
rect 11805 30141 11839 30175
rect 12448 30141 12482 30175
rect 12540 30141 12574 30175
rect 15577 30141 15611 30175
rect 16773 30141 16807 30175
rect 17325 30141 17359 30175
rect 18521 30141 18555 30175
rect 23949 30141 23983 30175
rect 26249 30141 26283 30175
rect 27629 30141 27663 30175
rect 30113 30141 30147 30175
rect 33333 30141 33367 30175
rect 34253 30141 34287 30175
rect 18245 30073 18279 30107
rect 20269 30073 20303 30107
rect 29285 30073 29319 30107
rect 31585 30073 31619 30107
rect 32413 30073 32447 30107
rect 36001 30073 36035 30107
rect 4813 30005 4847 30039
rect 5641 30005 5675 30039
rect 5825 30005 5859 30039
rect 10241 30005 10275 30039
rect 11713 30005 11747 30039
rect 13461 30005 13495 30039
rect 13645 30005 13679 30039
rect 14473 30005 14507 30039
rect 18705 30005 18739 30039
rect 24501 30005 24535 30039
rect 28733 30005 28767 30039
rect 33425 30005 33459 30039
rect 36553 30005 36587 30039
rect 37473 30005 37507 30039
rect 4445 29801 4479 29835
rect 12909 29801 12943 29835
rect 14749 29801 14783 29835
rect 23121 29801 23155 29835
rect 25513 29801 25547 29835
rect 26801 29801 26835 29835
rect 26985 29801 27019 29835
rect 27997 29801 28031 29835
rect 28457 29801 28491 29835
rect 28641 29801 28675 29835
rect 30113 29801 30147 29835
rect 32597 29801 32631 29835
rect 33885 29801 33919 29835
rect 12357 29733 12391 29767
rect 13369 29733 13403 29767
rect 14933 29733 14967 29767
rect 18245 29733 18279 29767
rect 31953 29733 31987 29767
rect 10701 29665 10735 29699
rect 14565 29665 14599 29699
rect 15945 29665 15979 29699
rect 18337 29665 18371 29699
rect 20821 29665 20855 29699
rect 31309 29665 31343 29699
rect 31493 29665 31527 29699
rect 36277 29665 36311 29699
rect 36461 29665 36495 29699
rect 38117 29665 38151 29699
rect 6193 29597 6227 29631
rect 7205 29597 7239 29631
rect 7297 29597 7331 29631
rect 7573 29597 7607 29631
rect 11345 29597 11379 29631
rect 11529 29597 11563 29631
rect 11805 29597 11839 29631
rect 12541 29597 12575 29631
rect 12633 29597 12667 29631
rect 13553 29597 13587 29631
rect 14473 29597 14507 29631
rect 14749 29597 14783 29631
rect 16221 29597 16255 29631
rect 17417 29597 17451 29631
rect 17969 29597 18003 29631
rect 18116 29597 18150 29631
rect 19257 29597 19291 29631
rect 19441 29597 19475 29631
rect 19625 29597 19659 29631
rect 23029 29597 23063 29631
rect 23673 29597 23707 29631
rect 24961 29597 24995 29631
rect 25513 29597 25547 29631
rect 25697 29597 25731 29631
rect 27445 29597 27479 29631
rect 27629 29597 27663 29631
rect 27813 29597 27847 29631
rect 30297 29597 30331 29631
rect 30389 29597 30423 29631
rect 30481 29597 30515 29631
rect 30757 29597 30791 29631
rect 33241 29597 33275 29631
rect 33425 29597 33459 29631
rect 34069 29597 34103 29631
rect 35541 29597 35575 29631
rect 5917 29529 5951 29563
rect 7389 29529 7423 29563
rect 10425 29529 10459 29563
rect 11161 29529 11195 29563
rect 11437 29529 11471 29563
rect 11667 29529 11701 29563
rect 19533 29529 19567 29563
rect 21097 29529 21131 29563
rect 26617 29529 26651 29563
rect 26833 29529 26867 29563
rect 27721 29529 27755 29563
rect 28825 29529 28859 29563
rect 30619 29529 30653 29563
rect 31585 29529 31619 29563
rect 32781 29529 32815 29563
rect 34713 29529 34747 29563
rect 34897 29529 34931 29563
rect 7021 29461 7055 29495
rect 8953 29461 8987 29495
rect 12725 29461 12759 29495
rect 17325 29461 17359 29495
rect 18613 29461 18647 29495
rect 19809 29461 19843 29495
rect 22569 29461 22603 29495
rect 23857 29461 23891 29495
rect 24869 29461 24903 29495
rect 28625 29461 28659 29495
rect 32413 29461 32447 29495
rect 32581 29461 32615 29495
rect 33333 29461 33367 29495
rect 35081 29461 35115 29495
rect 35633 29461 35667 29495
rect 7599 29257 7633 29291
rect 8585 29257 8619 29291
rect 10885 29257 10919 29291
rect 15945 29257 15979 29291
rect 18061 29257 18095 29291
rect 18429 29257 18463 29291
rect 20821 29257 20855 29291
rect 24317 29257 24351 29291
rect 26341 29257 26375 29291
rect 27353 29257 27387 29291
rect 28365 29257 28399 29291
rect 30941 29257 30975 29291
rect 32137 29257 32171 29291
rect 7389 29189 7423 29223
rect 12633 29189 12667 29223
rect 12817 29189 12851 29223
rect 14473 29189 14507 29223
rect 14565 29189 14599 29223
rect 15853 29189 15887 29223
rect 24225 29189 24259 29223
rect 25513 29189 25547 29223
rect 27261 29189 27295 29223
rect 31493 29189 31527 29223
rect 6561 29121 6595 29155
rect 8493 29121 8527 29155
rect 11805 29121 11839 29155
rect 12173 29121 12207 29155
rect 13645 29121 13679 29155
rect 13829 29121 13863 29155
rect 14289 29121 14323 29155
rect 14657 29121 14691 29155
rect 15761 29121 15795 29155
rect 16129 29121 16163 29155
rect 16681 29121 16715 29155
rect 16957 29121 16991 29155
rect 17325 29121 17359 29155
rect 18245 29121 18279 29155
rect 18337 29121 18371 29155
rect 19349 29121 19383 29155
rect 21005 29121 21039 29155
rect 21281 29121 21315 29155
rect 21833 29121 21867 29155
rect 26157 29121 26191 29155
rect 26433 29121 26467 29155
rect 27169 29121 27203 29155
rect 28549 29121 28583 29155
rect 28733 29121 28767 29155
rect 29101 29121 29135 29155
rect 29653 29121 29687 29155
rect 30389 29121 30423 29155
rect 30757 29121 30791 29155
rect 31401 29121 31435 29155
rect 31585 29121 31619 29155
rect 32137 29121 32171 29155
rect 32321 29121 32355 29155
rect 32965 29121 32999 29155
rect 33425 29121 33459 29155
rect 33885 29121 33919 29155
rect 34621 29121 34655 29155
rect 37565 29121 37599 29155
rect 6469 29053 6503 29087
rect 6929 29053 6963 29087
rect 9137 29053 9171 29087
rect 9413 29053 9447 29087
rect 11713 29053 11747 29087
rect 12081 29053 12115 29087
rect 13737 29053 13771 29087
rect 19073 29053 19107 29087
rect 22017 29053 22051 29087
rect 22293 29053 22327 29087
rect 25697 29053 25731 29087
rect 30297 29053 30331 29087
rect 33149 29053 33183 29087
rect 36369 29053 36403 29087
rect 11529 28985 11563 29019
rect 15577 28985 15611 29019
rect 18613 28985 18647 29019
rect 21189 28985 21223 29019
rect 26985 28985 27019 29019
rect 27537 28985 27571 29019
rect 32781 28985 32815 29019
rect 7573 28917 7607 28951
rect 7757 28917 7791 28951
rect 14841 28917 14875 28951
rect 17233 28917 17267 28951
rect 26157 28917 26191 28951
rect 30757 28917 30791 28951
rect 33333 28917 33367 28951
rect 33977 28917 34011 28951
rect 34878 28917 34912 28951
rect 37657 28917 37691 28951
rect 9137 28713 9171 28747
rect 11713 28713 11747 28747
rect 15853 28713 15887 28747
rect 19533 28713 19567 28747
rect 24409 28713 24443 28747
rect 28825 28713 28859 28747
rect 29009 28713 29043 28747
rect 30481 28713 30515 28747
rect 31585 28713 31619 28747
rect 34161 28713 34195 28747
rect 35541 28713 35575 28747
rect 9781 28645 9815 28679
rect 13093 28645 13127 28679
rect 18705 28645 18739 28679
rect 30021 28645 30055 28679
rect 7389 28577 7423 28611
rect 14105 28577 14139 28611
rect 16405 28577 16439 28611
rect 17325 28577 17359 28611
rect 17693 28577 17727 28611
rect 18429 28577 18463 28611
rect 21281 28577 21315 28611
rect 23581 28577 23615 28611
rect 26157 28577 26191 28611
rect 26801 28577 26835 28611
rect 33517 28577 33551 28611
rect 35081 28577 35115 28611
rect 37197 28577 37231 28611
rect 37933 28577 37967 28611
rect 7113 28509 7147 28543
rect 10793 28509 10827 28543
rect 11897 28509 11931 28543
rect 13001 28509 13035 28543
rect 13185 28509 13219 28543
rect 16497 28509 16531 28543
rect 16589 28509 16623 28543
rect 16681 28509 16715 28543
rect 17509 28509 17543 28543
rect 18337 28509 18371 28543
rect 21741 28509 21775 28543
rect 22569 28509 22603 28543
rect 23857 28509 23891 28543
rect 26893 28509 26927 28543
rect 26985 28509 27019 28543
rect 27077 28509 27111 28543
rect 27997 28509 28031 28543
rect 29561 28509 29595 28543
rect 29837 28509 29871 28543
rect 30665 28509 30699 28543
rect 30849 28509 30883 28543
rect 30941 28509 30975 28543
rect 31401 28509 31435 28543
rect 32321 28509 32355 28543
rect 33793 28509 33827 28543
rect 33977 28509 34011 28543
rect 34897 28509 34931 28543
rect 35541 28509 35575 28543
rect 35725 28509 35759 28543
rect 38117 28509 38151 28543
rect 9105 28441 9139 28475
rect 9321 28441 9355 28475
rect 9965 28441 9999 28475
rect 12081 28441 12115 28475
rect 14381 28441 14415 28475
rect 21005 28441 21039 28475
rect 22477 28441 22511 28475
rect 25881 28441 25915 28475
rect 27813 28441 27847 28475
rect 28641 28441 28675 28475
rect 28857 28441 28891 28475
rect 32413 28441 32447 28475
rect 32689 28441 32723 28475
rect 33675 28441 33709 28475
rect 33885 28441 33919 28475
rect 8953 28373 8987 28407
rect 10609 28373 10643 28407
rect 16865 28373 16899 28407
rect 21833 28373 21867 28407
rect 26617 28373 26651 28407
rect 27629 28373 27663 28407
rect 29653 28373 29687 28407
rect 32137 28373 32171 28407
rect 32505 28373 32539 28407
rect 34713 28373 34747 28407
rect 10241 28169 10275 28203
rect 14381 28169 14415 28203
rect 18429 28169 18463 28203
rect 20361 28169 20395 28203
rect 22017 28169 22051 28203
rect 22661 28169 22695 28203
rect 25881 28169 25915 28203
rect 26985 28169 27019 28203
rect 29745 28169 29779 28203
rect 32597 28169 32631 28203
rect 32765 28169 32799 28203
rect 36277 28169 36311 28203
rect 12817 28101 12851 28135
rect 15101 28101 15135 28135
rect 15301 28101 15335 28135
rect 15853 28101 15887 28135
rect 16957 28101 16991 28135
rect 21097 28101 21131 28135
rect 24869 28101 24903 28135
rect 27261 28101 27295 28135
rect 32965 28101 32999 28135
rect 33701 28101 33735 28135
rect 33793 28101 33827 28135
rect 34069 28101 34103 28135
rect 34805 28101 34839 28135
rect 6653 28033 6687 28067
rect 7757 28033 7791 28067
rect 8033 28033 8067 28067
rect 8217 28033 8251 28067
rect 9321 28033 9355 28067
rect 9413 28033 9447 28067
rect 10149 28033 10183 28067
rect 11713 28033 11747 28067
rect 12541 28033 12575 28067
rect 12725 28033 12759 28067
rect 12909 28033 12943 28067
rect 13553 28033 13587 28067
rect 14473 28033 14507 28067
rect 15945 28033 15979 28067
rect 16681 28033 16715 28067
rect 19073 28033 19107 28067
rect 19257 28033 19291 28067
rect 20177 28033 20211 28067
rect 20913 28033 20947 28067
rect 22109 28033 22143 28067
rect 22753 28033 22787 28067
rect 26065 28033 26099 28067
rect 26341 28033 26375 28067
rect 27169 28033 27203 28067
rect 27353 28033 27387 28067
rect 27537 28033 27571 28067
rect 28181 28033 28215 28067
rect 28917 28033 28951 28067
rect 29653 28033 29687 28067
rect 30389 28033 30423 28067
rect 31309 28033 31343 28067
rect 33563 28033 33597 28067
rect 33885 28033 33919 28067
rect 37841 28033 37875 28067
rect 9505 27965 9539 27999
rect 9597 27965 9631 27999
rect 11621 27965 11655 27999
rect 25145 27965 25179 27999
rect 26249 27965 26283 27999
rect 29101 27965 29135 27999
rect 33425 27965 33459 27999
rect 34529 27965 34563 27999
rect 12081 27897 12115 27931
rect 26157 27897 26191 27931
rect 28365 27897 28399 27931
rect 6561 27829 6595 27863
rect 7573 27829 7607 27863
rect 9137 27829 9171 27863
rect 13093 27829 13127 27863
rect 13737 27829 13771 27863
rect 14933 27829 14967 27863
rect 15117 27829 15151 27863
rect 18889 27829 18923 27863
rect 23397 27829 23431 27863
rect 30481 27829 30515 27863
rect 31493 27829 31527 27863
rect 32781 27829 32815 27863
rect 6579 27625 6613 27659
rect 7297 27625 7331 27659
rect 11805 27625 11839 27659
rect 13289 27625 13323 27659
rect 16681 27625 16715 27659
rect 17601 27625 17635 27659
rect 19257 27625 19291 27659
rect 28365 27625 28399 27659
rect 33977 27625 34011 27659
rect 18061 27557 18095 27591
rect 23765 27557 23799 27591
rect 24501 27557 24535 27591
rect 28641 27557 28675 27591
rect 34713 27557 34747 27591
rect 6837 27489 6871 27523
rect 9597 27489 9631 27523
rect 9689 27489 9723 27523
rect 10977 27489 11011 27523
rect 17693 27489 17727 27523
rect 19625 27489 19659 27523
rect 20269 27489 20303 27523
rect 25605 27489 25639 27523
rect 26433 27489 26467 27523
rect 26525 27489 26559 27523
rect 31309 27489 31343 27523
rect 31493 27489 31527 27523
rect 32321 27489 32355 27523
rect 38117 27489 38151 27523
rect 7481 27421 7515 27455
rect 7849 27421 7883 27455
rect 9505 27421 9539 27455
rect 9781 27421 9815 27455
rect 10885 27421 10919 27455
rect 11069 27421 11103 27455
rect 13553 27421 13587 27455
rect 14289 27421 14323 27455
rect 14933 27421 14967 27455
rect 15485 27421 15519 27455
rect 15577 27421 15611 27455
rect 16221 27421 16255 27455
rect 16313 27421 16347 27455
rect 16497 27421 16531 27455
rect 17877 27421 17911 27455
rect 18521 27421 18555 27455
rect 19441 27421 19475 27455
rect 19717 27421 19751 27455
rect 20177 27421 20211 27455
rect 20361 27421 20395 27455
rect 21005 27421 21039 27455
rect 22661 27421 22695 27455
rect 23673 27421 23707 27455
rect 24685 27421 24719 27455
rect 25697 27421 25731 27455
rect 26341 27421 26375 27455
rect 26617 27421 26651 27455
rect 27169 27421 27203 27455
rect 27353 27421 27387 27455
rect 27537 27421 27571 27455
rect 28365 27421 28399 27455
rect 28457 27421 28491 27455
rect 29561 27421 29595 27455
rect 30205 27421 30239 27455
rect 30481 27421 30515 27455
rect 31217 27421 31251 27455
rect 31401 27421 31435 27455
rect 32597 27421 32631 27455
rect 34897 27421 34931 27455
rect 35173 27421 35207 27455
rect 36277 27421 36311 27455
rect 7573 27353 7607 27387
rect 7665 27353 7699 27387
rect 14841 27353 14875 27387
rect 17601 27353 17635 27387
rect 27445 27353 27479 27387
rect 28181 27353 28215 27387
rect 30297 27353 30331 27387
rect 33793 27353 33827 27387
rect 35081 27353 35115 27387
rect 36461 27353 36495 27387
rect 5089 27285 5123 27319
rect 9321 27285 9355 27319
rect 14105 27285 14139 27319
rect 15761 27285 15795 27319
rect 18613 27285 18647 27319
rect 20913 27285 20947 27319
rect 22753 27285 22787 27319
rect 26157 27285 26191 27319
rect 27721 27285 27755 27319
rect 29653 27285 29687 27319
rect 30665 27285 30699 27319
rect 31677 27285 31711 27319
rect 33993 27285 34027 27319
rect 34161 27285 34195 27319
rect 8861 27081 8895 27115
rect 11713 27081 11747 27115
rect 18705 27081 18739 27115
rect 18889 27081 18923 27115
rect 21081 27081 21115 27115
rect 28825 27081 28859 27115
rect 31309 27081 31343 27115
rect 31585 27081 31619 27115
rect 32965 27081 32999 27115
rect 34713 27081 34747 27115
rect 37381 27081 37415 27115
rect 21281 27013 21315 27047
rect 24409 27013 24443 27047
rect 29837 27013 29871 27047
rect 29975 27013 30009 27047
rect 31401 27013 31435 27047
rect 33977 27013 34011 27047
rect 34161 27013 34195 27047
rect 6469 26945 6503 26979
rect 11897 26945 11931 26979
rect 15669 26945 15703 26979
rect 15853 26945 15887 26979
rect 15945 26945 15979 26979
rect 16865 26945 16899 26979
rect 16957 26945 16991 26979
rect 17877 26945 17911 26979
rect 18797 26945 18831 26979
rect 19073 26945 19107 26979
rect 19717 26945 19751 26979
rect 19901 26945 19935 26979
rect 21833 26945 21867 26979
rect 29653 26945 29687 26979
rect 29745 26945 29779 26979
rect 31217 26945 31251 26979
rect 32321 26945 32355 26979
rect 33149 26945 33183 26979
rect 33425 26945 33459 26979
rect 34621 26945 34655 26979
rect 35265 26945 35299 26979
rect 35449 26945 35483 26979
rect 37473 26945 37507 26979
rect 6745 26877 6779 26911
rect 8217 26877 8251 26911
rect 10333 26877 10367 26911
rect 10609 26877 10643 26911
rect 13277 26877 13311 26911
rect 13553 26877 13587 26911
rect 15025 26877 15059 26911
rect 17693 26877 17727 26911
rect 19533 26877 19567 26911
rect 19809 26877 19843 26911
rect 19993 26877 20027 26911
rect 22109 26877 22143 26911
rect 24133 26877 24167 26911
rect 27077 26877 27111 26911
rect 27353 26877 27387 26911
rect 30113 26877 30147 26911
rect 33333 26877 33367 26911
rect 23581 26809 23615 26843
rect 31033 26809 31067 26843
rect 15485 26741 15519 26775
rect 16681 26741 16715 26775
rect 18061 26741 18095 26775
rect 18521 26741 18555 26775
rect 20913 26741 20947 26775
rect 21097 26741 21131 26775
rect 25881 26741 25915 26775
rect 29469 26741 29503 26775
rect 32413 26741 32447 26775
rect 33425 26741 33459 26775
rect 35265 26741 35299 26775
rect 7021 26537 7055 26571
rect 10425 26537 10459 26571
rect 24777 26537 24811 26571
rect 25881 26537 25915 26571
rect 26801 26537 26835 26571
rect 31953 26537 31987 26571
rect 34713 26537 34747 26571
rect 7665 26469 7699 26503
rect 15577 26469 15611 26503
rect 16957 26469 16991 26503
rect 19349 26469 19383 26503
rect 22293 26469 22327 26503
rect 26249 26469 26283 26503
rect 28273 26469 28307 26503
rect 31217 26469 31251 26503
rect 34161 26469 34195 26503
rect 8217 26401 8251 26435
rect 8953 26401 8987 26435
rect 9873 26401 9907 26435
rect 14749 26401 14783 26435
rect 16129 26401 16163 26435
rect 18521 26401 18555 26435
rect 21097 26401 21131 26435
rect 25973 26401 26007 26435
rect 27077 26401 27111 26435
rect 27261 26401 27295 26435
rect 28733 26401 28767 26435
rect 28917 26401 28951 26435
rect 30113 26401 30147 26435
rect 32597 26401 32631 26435
rect 1961 26333 1995 26367
rect 7205 26333 7239 26367
rect 8125 26333 8159 26367
rect 9137 26333 9171 26367
rect 9781 26333 9815 26367
rect 9965 26333 9999 26367
rect 10609 26333 10643 26367
rect 11989 26333 12023 26367
rect 12173 26333 12207 26367
rect 14105 26333 14139 26367
rect 14933 26333 14967 26367
rect 15117 26333 15151 26367
rect 15945 26333 15979 26367
rect 17141 26333 17175 26367
rect 18337 26333 18371 26367
rect 18429 26333 18463 26367
rect 21741 26333 21775 26367
rect 22569 26333 22603 26367
rect 22845 26333 22879 26367
rect 23397 26333 23431 26367
rect 23673 26333 23707 26367
rect 24593 26333 24627 26367
rect 25789 26333 25823 26367
rect 26065 26333 26099 26367
rect 26985 26333 27019 26367
rect 27169 26333 27203 26367
rect 28641 26333 28675 26367
rect 30271 26333 30305 26367
rect 30572 26333 30606 26367
rect 31401 26333 31435 26367
rect 32137 26333 32171 26367
rect 32321 26333 32355 26367
rect 33609 26333 33643 26367
rect 33793 26333 33827 26367
rect 33977 26333 34011 26367
rect 34897 26333 34931 26367
rect 34989 26333 35023 26367
rect 35541 26333 35575 26367
rect 35725 26333 35759 26367
rect 37013 26333 37047 26367
rect 37841 26333 37875 26367
rect 8033 26265 8067 26299
rect 16037 26265 16071 26299
rect 20821 26265 20855 26299
rect 24409 26265 24443 26299
rect 30389 26265 30423 26299
rect 30481 26265 30515 26299
rect 32229 26265 32263 26299
rect 32459 26265 32493 26299
rect 33885 26265 33919 26299
rect 35633 26265 35667 26299
rect 9321 26197 9355 26231
rect 12081 26197 12115 26231
rect 14289 26197 14323 26231
rect 17969 26197 18003 26231
rect 21557 26197 21591 26231
rect 30757 26197 30791 26231
rect 7389 25993 7423 26027
rect 10149 25993 10183 26027
rect 14289 25993 14323 26027
rect 15577 25993 15611 26027
rect 18429 25993 18463 26027
rect 22109 25993 22143 26027
rect 22477 25993 22511 26027
rect 24869 25993 24903 26027
rect 27353 25993 27387 26027
rect 27905 25993 27939 26027
rect 33425 25993 33459 26027
rect 36093 25993 36127 26027
rect 9413 25925 9447 25959
rect 11980 25925 12014 25959
rect 16957 25925 16991 25959
rect 21081 25925 21115 25959
rect 21281 25925 21315 25959
rect 26433 25925 26467 25959
rect 26985 25925 27019 25959
rect 27185 25925 27219 25959
rect 28089 25925 28123 25959
rect 33793 25925 33827 25959
rect 34621 25925 34655 25959
rect 1869 25857 1903 25891
rect 7297 25857 7331 25891
rect 9321 25857 9355 25891
rect 9597 25857 9631 25891
rect 10241 25857 10275 25891
rect 11713 25857 11747 25891
rect 14197 25857 14231 25891
rect 15117 25857 15151 25891
rect 15853 25857 15887 25891
rect 16681 25857 16715 25891
rect 19441 25857 19475 25891
rect 20453 25857 20487 25891
rect 22293 25857 22327 25891
rect 22569 25857 22603 25891
rect 23121 25857 23155 25891
rect 23305 25857 23339 25891
rect 23489 25857 23523 25891
rect 23581 25857 23615 25891
rect 24133 25857 24167 25891
rect 24777 25857 24811 25891
rect 25421 25857 25455 25891
rect 25605 25857 25639 25891
rect 26249 25857 26283 25891
rect 27813 25857 27847 25891
rect 28825 25857 28859 25891
rect 29929 25857 29963 25891
rect 30205 25857 30239 25891
rect 30665 25857 30699 25891
rect 32413 25857 32447 25891
rect 33609 25857 33643 25891
rect 33885 25857 33919 25891
rect 34345 25857 34379 25891
rect 37289 25857 37323 25891
rect 2053 25789 2087 25823
rect 2881 25789 2915 25823
rect 15577 25789 15611 25823
rect 15761 25789 15795 25823
rect 28641 25789 28675 25823
rect 30941 25789 30975 25823
rect 32137 25789 32171 25823
rect 19625 25721 19659 25755
rect 20913 25721 20947 25755
rect 24317 25721 24351 25755
rect 28089 25721 28123 25755
rect 9597 25653 9631 25687
rect 13093 25653 13127 25687
rect 15025 25653 15059 25687
rect 20269 25653 20303 25687
rect 21097 25653 21131 25687
rect 25513 25653 25547 25687
rect 26065 25653 26099 25687
rect 27169 25653 27203 25687
rect 37381 25653 37415 25687
rect 38117 25653 38151 25687
rect 2789 25449 2823 25483
rect 11805 25449 11839 25483
rect 16129 25449 16163 25483
rect 17417 25449 17451 25483
rect 19441 25449 19475 25483
rect 22385 25449 22419 25483
rect 24501 25449 24535 25483
rect 25513 25449 25547 25483
rect 27537 25449 27571 25483
rect 29745 25449 29779 25483
rect 32045 25449 32079 25483
rect 32781 25449 32815 25483
rect 35449 25449 35483 25483
rect 20269 25381 20303 25415
rect 33425 25381 33459 25415
rect 34713 25381 34747 25415
rect 6653 25313 6687 25347
rect 9597 25313 9631 25347
rect 14105 25313 14139 25347
rect 21281 25313 21315 25347
rect 30573 25313 30607 25347
rect 36277 25313 36311 25347
rect 36461 25313 36495 25347
rect 38117 25313 38151 25347
rect 2881 25245 2915 25279
rect 9137 25245 9171 25279
rect 12081 25245 12115 25279
rect 12173 25245 12207 25279
rect 12265 25245 12299 25279
rect 12449 25245 12483 25279
rect 13461 25245 13495 25279
rect 17325 25245 17359 25279
rect 18061 25245 18095 25279
rect 19257 25245 19291 25279
rect 20913 25245 20947 25279
rect 22569 25245 22603 25279
rect 22753 25245 22787 25279
rect 23305 25245 23339 25279
rect 23489 25245 23523 25279
rect 24685 25245 24719 25279
rect 25697 25245 25731 25279
rect 25973 25245 26007 25279
rect 26617 25245 26651 25279
rect 26893 25245 26927 25279
rect 28273 25245 28307 25279
rect 29653 25245 29687 25279
rect 29837 25245 29871 25279
rect 30297 25245 30331 25279
rect 32873 25245 32907 25279
rect 33333 25245 33367 25279
rect 33609 25245 33643 25279
rect 34713 25245 34747 25279
rect 34897 25245 34931 25279
rect 35357 25245 35391 25279
rect 6920 25177 6954 25211
rect 9864 25177 9898 25211
rect 14372 25177 14406 25211
rect 16313 25177 16347 25211
rect 20085 25177 20119 25211
rect 25881 25177 25915 25211
rect 27521 25177 27555 25211
rect 27721 25177 27755 25211
rect 8033 25109 8067 25143
rect 9045 25109 9079 25143
rect 10977 25109 11011 25143
rect 13369 25109 13403 25143
rect 15485 25109 15519 25143
rect 15945 25109 15979 25143
rect 16113 25109 16147 25143
rect 18245 25109 18279 25143
rect 26433 25109 26467 25143
rect 26801 25109 26835 25143
rect 27353 25109 27387 25143
rect 28365 25109 28399 25143
rect 33793 25109 33827 25143
rect 8677 24905 8711 24939
rect 12081 24905 12115 24939
rect 14749 24905 14783 24939
rect 15117 24905 15151 24939
rect 25881 24905 25915 24939
rect 29469 24905 29503 24939
rect 8309 24837 8343 24871
rect 8509 24837 8543 24871
rect 19165 24837 19199 24871
rect 20361 24837 20395 24871
rect 6837 24769 6871 24803
rect 7021 24769 7055 24803
rect 7665 24769 7699 24803
rect 7849 24769 7883 24803
rect 9781 24769 9815 24803
rect 9873 24769 9907 24803
rect 9965 24769 9999 24803
rect 10149 24769 10183 24803
rect 11897 24769 11931 24803
rect 12173 24769 12207 24803
rect 12817 24769 12851 24803
rect 13461 24769 13495 24803
rect 13645 24769 13679 24803
rect 14289 24769 14323 24803
rect 14933 24769 14967 24803
rect 15209 24769 15243 24803
rect 15945 24769 15979 24803
rect 17049 24769 17083 24803
rect 17141 24769 17175 24803
rect 21189 24769 21223 24803
rect 21833 24769 21867 24803
rect 25973 24769 26007 24803
rect 27169 24769 27203 24803
rect 30021 24769 30055 24803
rect 30205 24769 30239 24803
rect 30389 24769 30423 24803
rect 30849 24769 30883 24803
rect 30941 24769 30975 24803
rect 31125 24769 31159 24803
rect 34345 24769 34379 24803
rect 7481 24701 7515 24735
rect 13553 24701 13587 24735
rect 15669 24701 15703 24735
rect 15761 24701 15795 24735
rect 17693 24701 17727 24735
rect 19441 24701 19475 24735
rect 22109 24701 22143 24735
rect 23305 24701 23339 24735
rect 23581 24701 23615 24735
rect 25053 24701 25087 24735
rect 26157 24701 26191 24735
rect 27721 24701 27755 24735
rect 27997 24701 28031 24735
rect 32137 24701 32171 24735
rect 32413 24701 32447 24735
rect 33885 24701 33919 24735
rect 34621 24701 34655 24735
rect 36093 24701 36127 24735
rect 12725 24633 12759 24667
rect 30849 24633 30883 24667
rect 6929 24565 6963 24599
rect 8493 24565 8527 24599
rect 9505 24565 9539 24599
rect 11897 24565 11931 24599
rect 14197 24565 14231 24599
rect 16129 24565 16163 24599
rect 25513 24565 25547 24599
rect 26985 24565 27019 24599
rect 36553 24565 36587 24599
rect 37841 24565 37875 24599
rect 7573 24361 7607 24395
rect 9137 24361 9171 24395
rect 9873 24361 9907 24395
rect 13093 24361 13127 24395
rect 14933 24361 14967 24395
rect 15117 24361 15151 24395
rect 18613 24361 18647 24395
rect 24409 24361 24443 24395
rect 25697 24361 25731 24395
rect 27905 24361 27939 24395
rect 28365 24361 28399 24395
rect 32505 24361 32539 24395
rect 33149 24361 33183 24395
rect 34805 24361 34839 24395
rect 13277 24293 13311 24327
rect 14197 24293 14231 24327
rect 17877 24293 17911 24327
rect 20453 24293 20487 24327
rect 23765 24293 23799 24327
rect 8953 24225 8987 24259
rect 15485 24225 15519 24259
rect 21557 24225 21591 24259
rect 26433 24225 26467 24259
rect 29561 24225 29595 24259
rect 36277 24225 36311 24259
rect 7021 24157 7055 24191
rect 7757 24157 7791 24191
rect 7849 24157 7883 24191
rect 8217 24157 8251 24191
rect 9229 24157 9263 24191
rect 9689 24157 9723 24191
rect 9873 24157 9907 24191
rect 10609 24157 10643 24191
rect 17325 24157 17359 24191
rect 17969 24157 18003 24191
rect 18429 24157 18463 24191
rect 19257 24157 19291 24191
rect 21833 24157 21867 24191
rect 22477 24157 22511 24191
rect 23673 24157 23707 24191
rect 24593 24157 24627 24191
rect 25421 24157 25455 24191
rect 25513 24157 25547 24191
rect 26157 24157 26191 24191
rect 28549 24157 28583 24191
rect 31953 24157 31987 24191
rect 32597 24157 32631 24191
rect 33057 24157 33091 24191
rect 34161 24157 34195 24191
rect 34713 24157 34747 24191
rect 35541 24157 35575 24191
rect 6837 24089 6871 24123
rect 7941 24089 7975 24123
rect 8079 24089 8113 24123
rect 10876 24089 10910 24123
rect 12909 24089 12943 24123
rect 13109 24089 13143 24123
rect 14381 24089 14415 24123
rect 15117 24089 15151 24123
rect 17058 24089 17092 24123
rect 19441 24089 19475 24123
rect 20269 24089 20303 24123
rect 23029 24089 23063 24123
rect 29837 24089 29871 24123
rect 31861 24089 31895 24123
rect 36461 24089 36495 24123
rect 38117 24089 38151 24123
rect 6653 24021 6687 24055
rect 8953 24021 8987 24055
rect 11989 24021 12023 24055
rect 15945 24021 15979 24055
rect 31309 24021 31343 24055
rect 35449 24021 35483 24055
rect 7665 23817 7699 23851
rect 10241 23817 10275 23851
rect 11529 23817 11563 23851
rect 15117 23817 15151 23851
rect 19993 23817 20027 23851
rect 24133 23817 24167 23851
rect 24501 23817 24535 23851
rect 25421 23817 25455 23851
rect 27353 23817 27387 23851
rect 37381 23817 37415 23851
rect 6745 23749 6779 23783
rect 15485 23749 15519 23783
rect 26157 23749 26191 23783
rect 6561 23681 6595 23715
rect 6653 23681 6687 23715
rect 6863 23681 6897 23715
rect 7849 23681 7883 23715
rect 7941 23681 7975 23715
rect 8125 23681 8159 23715
rect 8861 23681 8895 23715
rect 9597 23681 9631 23715
rect 9781 23681 9815 23715
rect 10425 23681 10459 23715
rect 11713 23681 11747 23715
rect 11805 23681 11839 23715
rect 11897 23681 11931 23715
rect 12015 23681 12049 23715
rect 12173 23681 12207 23715
rect 12817 23681 12851 23715
rect 13073 23681 13107 23715
rect 15320 23681 15354 23715
rect 15577 23681 15611 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 18438 23681 18472 23715
rect 18705 23681 18739 23715
rect 19625 23681 19659 23715
rect 19809 23681 19843 23715
rect 20545 23681 20579 23715
rect 20729 23681 20763 23715
rect 21833 23681 21867 23715
rect 24317 23681 24351 23715
rect 24593 23681 24627 23715
rect 25421 23681 25455 23715
rect 26249 23681 26283 23715
rect 27445 23681 27479 23715
rect 30757 23681 30791 23715
rect 32873 23681 32907 23715
rect 33517 23681 33551 23715
rect 33977 23681 34011 23715
rect 36277 23681 36311 23715
rect 37289 23681 37323 23715
rect 37933 23681 37967 23715
rect 7021 23613 7055 23647
rect 8033 23613 8067 23647
rect 16773 23613 16807 23647
rect 20453 23613 20487 23647
rect 22109 23613 22143 23647
rect 25053 23613 25087 23647
rect 25605 23613 25639 23647
rect 34253 23613 34287 23647
rect 8677 23545 8711 23579
rect 14197 23545 14231 23579
rect 30941 23545 30975 23579
rect 6377 23477 6411 23511
rect 9413 23477 9447 23511
rect 17325 23477 17359 23511
rect 23581 23477 23615 23511
rect 33425 23477 33459 23511
rect 35725 23477 35759 23511
rect 36369 23477 36403 23511
rect 38025 23477 38059 23511
rect 6653 23273 6687 23307
rect 10333 23273 10367 23307
rect 11253 23273 11287 23307
rect 12909 23273 12943 23307
rect 15485 23273 15519 23307
rect 16865 23273 16899 23307
rect 21465 23273 21499 23307
rect 22017 23273 22051 23307
rect 35449 23273 35483 23307
rect 21373 23205 21407 23239
rect 7757 23137 7791 23171
rect 11161 23137 11195 23171
rect 15025 23137 15059 23171
rect 15577 23137 15611 23171
rect 19993 23137 20027 23171
rect 22201 23137 22235 23171
rect 22293 23137 22327 23171
rect 22385 23137 22419 23171
rect 29561 23137 29595 23171
rect 32045 23137 32079 23171
rect 36369 23137 36403 23171
rect 38025 23137 38059 23171
rect 5273 23069 5307 23103
rect 5540 23069 5574 23103
rect 7481 23069 7515 23103
rect 8953 23069 8987 23103
rect 10793 23069 10827 23103
rect 11253 23069 11287 23103
rect 12081 23069 12115 23103
rect 12173 23069 12207 23103
rect 13093 23069 13127 23103
rect 13277 23069 13311 23103
rect 13395 23069 13429 23103
rect 13553 23069 13587 23103
rect 14657 23069 14691 23103
rect 15761 23069 15795 23103
rect 17141 23069 17175 23103
rect 17233 23069 17267 23103
rect 17325 23069 17359 23103
rect 17509 23069 17543 23103
rect 17969 23069 18003 23103
rect 18153 23069 18187 23103
rect 19533 23069 19567 23103
rect 19809 23069 19843 23103
rect 20637 23069 20671 23103
rect 21189 23069 21223 23103
rect 21281 23069 21315 23103
rect 21557 23069 21591 23103
rect 22477 23069 22511 23103
rect 23673 23069 23707 23103
rect 25605 23069 25639 23103
rect 26433 23069 26467 23103
rect 27077 23069 27111 23103
rect 27721 23069 27755 23103
rect 35265 23069 35299 23103
rect 36185 23069 36219 23103
rect 9198 23001 9232 23035
rect 11897 23001 11931 23035
rect 13185 23001 13219 23035
rect 14749 23001 14783 23035
rect 15485 23001 15519 23035
rect 23857 23001 23891 23035
rect 24409 23001 24443 23035
rect 24593 23001 24627 23035
rect 24961 23001 24995 23035
rect 29837 23001 29871 23035
rect 32321 23001 32355 23035
rect 11437 22933 11471 22967
rect 12265 22933 12299 22967
rect 12449 22933 12483 22967
rect 14473 22933 14507 22967
rect 14841 22933 14875 22967
rect 15945 22933 15979 22967
rect 18061 22933 18095 22967
rect 19625 22933 19659 22967
rect 20545 22933 20579 22967
rect 23489 22933 23523 22967
rect 24685 22933 24719 22967
rect 24777 22933 24811 22967
rect 25513 22933 25547 22967
rect 26525 22933 26559 22967
rect 27261 22933 27295 22967
rect 27813 22933 27847 22967
rect 31309 22933 31343 22967
rect 33793 22933 33827 22967
rect 8769 22729 8803 22763
rect 9505 22729 9539 22763
rect 10609 22729 10643 22763
rect 11897 22729 11931 22763
rect 12081 22729 12115 22763
rect 12541 22729 12575 22763
rect 13553 22729 13587 22763
rect 17141 22729 17175 22763
rect 18981 22729 19015 22763
rect 19625 22729 19659 22763
rect 29469 22729 29503 22763
rect 33517 22729 33551 22763
rect 6745 22661 6779 22695
rect 7573 22661 7607 22695
rect 9597 22661 9631 22695
rect 9781 22661 9815 22695
rect 13921 22661 13955 22695
rect 14473 22661 14507 22695
rect 18889 22661 18923 22695
rect 27261 22661 27295 22695
rect 4353 22593 4387 22627
rect 4620 22593 4654 22627
rect 6377 22593 6411 22627
rect 6561 22593 6595 22627
rect 6653 22593 6687 22627
rect 6863 22593 6897 22627
rect 7665 22593 7699 22627
rect 8217 22593 8251 22627
rect 8493 22593 8527 22627
rect 8585 22593 8619 22627
rect 9413 22593 9447 22627
rect 10425 22593 10459 22627
rect 10701 22593 10735 22627
rect 10793 22593 10827 22627
rect 11713 22593 11747 22627
rect 11805 22593 11839 22627
rect 13001 22593 13035 22627
rect 13737 22593 13771 22627
rect 14013 22593 14047 22627
rect 14657 22593 14691 22627
rect 15393 22593 15427 22627
rect 15669 22593 15703 22627
rect 15853 22593 15887 22627
rect 16129 22593 16163 22627
rect 16957 22593 16991 22627
rect 17233 22593 17267 22627
rect 18153 22593 18187 22627
rect 18705 22593 18739 22627
rect 18981 22593 19015 22627
rect 20821 22593 20855 22627
rect 21097 22593 21131 22627
rect 26157 22593 26191 22627
rect 29285 22593 29319 22627
rect 30113 22593 30147 22627
rect 30573 22593 30607 22627
rect 32321 22593 32355 22627
rect 32965 22593 32999 22627
rect 33425 22593 33459 22627
rect 34437 22593 34471 22627
rect 34897 22593 34931 22627
rect 37289 22593 37323 22627
rect 37933 22593 37967 22627
rect 7021 22525 7055 22559
rect 11529 22525 11563 22559
rect 12725 22525 12759 22559
rect 12817 22525 12851 22559
rect 12909 22525 12943 22559
rect 15301 22525 15335 22559
rect 19993 22525 20027 22559
rect 22477 22525 22511 22559
rect 22753 22525 22787 22559
rect 23765 22525 23799 22559
rect 24041 22525 24075 22559
rect 26985 22525 27019 22559
rect 34161 22525 34195 22559
rect 35081 22525 35115 22559
rect 36737 22525 36771 22559
rect 9229 22457 9263 22491
rect 16957 22457 16991 22491
rect 20821 22457 20855 22491
rect 25973 22457 26007 22491
rect 32873 22457 32907 22491
rect 34345 22457 34379 22491
rect 38025 22457 38059 22491
rect 5733 22389 5767 22423
rect 8309 22389 8343 22423
rect 10701 22389 10735 22423
rect 18061 22389 18095 22423
rect 19441 22389 19475 22423
rect 19625 22389 19659 22423
rect 25513 22389 25547 22423
rect 28733 22389 28767 22423
rect 30021 22389 30055 22423
rect 30757 22389 30791 22423
rect 32229 22389 32263 22423
rect 34437 22389 34471 22423
rect 37381 22389 37415 22423
rect 6653 22185 6687 22219
rect 9137 22185 9171 22219
rect 10425 22185 10459 22219
rect 15393 22185 15427 22219
rect 17693 22185 17727 22219
rect 20453 22185 20487 22219
rect 25053 22185 25087 22219
rect 33057 22185 33091 22219
rect 33793 22185 33827 22219
rect 33977 22185 34011 22219
rect 35357 22185 35391 22219
rect 7481 22117 7515 22151
rect 11207 22117 11241 22151
rect 12265 22049 12299 22083
rect 14105 22049 14139 22083
rect 15761 22049 15795 22083
rect 16957 22049 16991 22083
rect 19901 22049 19935 22083
rect 20269 22049 20303 22083
rect 22017 22049 22051 22083
rect 25789 22049 25823 22083
rect 27537 22049 27571 22083
rect 30481 22049 30515 22083
rect 32873 22049 32907 22083
rect 37473 22049 37507 22083
rect 37933 22049 37967 22083
rect 38117 22049 38151 22083
rect 6377 21981 6411 22015
rect 6653 21981 6687 22015
rect 7021 21981 7055 22015
rect 7665 21981 7699 22015
rect 7849 21981 7883 22015
rect 8953 21981 8987 22015
rect 9137 21981 9171 22015
rect 10609 21981 10643 22015
rect 11069 21981 11103 22015
rect 11345 21981 11379 22015
rect 11529 21981 11563 22015
rect 12541 21981 12575 22015
rect 14381 21981 14415 22015
rect 15577 21981 15611 22015
rect 16313 21981 16347 22015
rect 16497 21981 16531 22015
rect 16589 21981 16623 22015
rect 16681 21981 16715 22015
rect 17417 21981 17451 22015
rect 18613 21981 18647 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 22293 21981 22327 22015
rect 22937 21981 22971 22015
rect 23581 21981 23615 22015
rect 23765 21981 23799 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 28181 21981 28215 22015
rect 28365 21981 28399 22015
rect 29009 21981 29043 22015
rect 30021 21981 30055 22015
rect 33057 21981 33091 22015
rect 35081 21981 35115 22015
rect 35173 21981 35207 22015
rect 8033 21913 8067 21947
rect 17693 21913 17727 21947
rect 18429 21913 18463 21947
rect 22753 21913 22787 21947
rect 23121 21913 23155 21947
rect 26065 21913 26099 21947
rect 29929 21913 29963 21947
rect 30757 21913 30791 21947
rect 32781 21913 32815 21947
rect 34161 21913 34195 21947
rect 35357 21913 35391 21947
rect 6837 21845 6871 21879
rect 7757 21845 7791 21879
rect 11529 21845 11563 21879
rect 17509 21845 17543 21879
rect 19257 21845 19291 21879
rect 20085 21845 20119 21879
rect 23765 21845 23799 21879
rect 24409 21845 24443 21879
rect 28181 21845 28215 21879
rect 28917 21845 28951 21879
rect 32229 21845 32263 21879
rect 33241 21845 33275 21879
rect 33961 21845 33995 21879
rect 34897 21845 34931 21879
rect 5733 21641 5767 21675
rect 10517 21641 10551 21675
rect 12909 21641 12943 21675
rect 23581 21641 23615 21675
rect 30757 21641 30791 21675
rect 7665 21573 7699 21607
rect 7941 21573 7975 21607
rect 8033 21573 8067 21607
rect 8171 21573 8205 21607
rect 17816 21573 17850 21607
rect 18705 21573 18739 21607
rect 19625 21573 19659 21607
rect 25239 21573 25273 21607
rect 26985 21573 27019 21607
rect 32873 21573 32907 21607
rect 35081 21573 35115 21607
rect 4353 21505 4387 21539
rect 4620 21505 4654 21539
rect 6377 21505 6411 21539
rect 7849 21505 7883 21539
rect 9404 21505 9438 21539
rect 11529 21505 11563 21539
rect 11785 21505 11819 21539
rect 13553 21505 13587 21539
rect 13737 21505 13771 21539
rect 13921 21505 13955 21539
rect 14381 21505 14415 21539
rect 14565 21505 14599 21539
rect 15945 21505 15979 21539
rect 19349 21505 19383 21539
rect 19441 21505 19475 21539
rect 20269 21505 20303 21539
rect 20453 21505 20487 21539
rect 21097 21505 21131 21539
rect 21833 21505 21867 21539
rect 22109 21505 22143 21539
rect 23397 21505 23431 21539
rect 23673 21505 23707 21539
rect 24593 21505 24627 21539
rect 26341 21505 26375 21539
rect 26433 21505 26467 21539
rect 27169 21505 27203 21539
rect 27261 21505 27295 21539
rect 30665 21505 30699 21539
rect 30849 21505 30883 21539
rect 32137 21505 32171 21539
rect 32321 21505 32355 21539
rect 32965 21505 32999 21539
rect 33241 21505 33275 21539
rect 33425 21505 33459 21539
rect 33701 21505 33735 21539
rect 34161 21505 34195 21539
rect 37657 21505 37691 21539
rect 6653 21437 6687 21471
rect 8309 21437 8343 21471
rect 9137 21437 9171 21471
rect 15761 21437 15795 21471
rect 18061 21437 18095 21471
rect 20913 21437 20947 21471
rect 26157 21437 26191 21471
rect 28273 21437 28307 21471
rect 28549 21437 28583 21471
rect 34805 21437 34839 21471
rect 16129 21369 16163 21403
rect 19625 21369 19659 21403
rect 25421 21369 25455 21403
rect 26433 21369 26467 21403
rect 26985 21369 27019 21403
rect 30481 21369 30515 21403
rect 14749 21301 14783 21335
rect 16681 21301 16715 21335
rect 18613 21301 18647 21335
rect 20361 21301 20395 21335
rect 21281 21301 21315 21335
rect 23397 21301 23431 21335
rect 24501 21301 24535 21335
rect 30021 21301 30055 21335
rect 31033 21301 31067 21335
rect 32229 21301 32263 21335
rect 34253 21301 34287 21335
rect 36553 21301 36587 21335
rect 37749 21301 37783 21335
rect 5365 21097 5399 21131
rect 6377 21097 6411 21131
rect 8217 21097 8251 21131
rect 10517 21097 10551 21131
rect 13369 21097 13403 21131
rect 21189 21097 21223 21131
rect 25899 21097 25933 21131
rect 26617 21097 26651 21131
rect 27905 21097 27939 21131
rect 28365 21097 28399 21131
rect 30021 21097 30055 21131
rect 30297 21097 30331 21131
rect 33701 21097 33735 21131
rect 34069 21097 34103 21131
rect 9413 21029 9447 21063
rect 27169 21029 27203 21063
rect 30941 21029 30975 21063
rect 35633 21029 35667 21063
rect 5917 20961 5951 20995
rect 6193 20961 6227 20995
rect 11161 20961 11195 20995
rect 11621 20961 11655 20995
rect 12817 20961 12851 20995
rect 16773 20961 16807 20995
rect 18521 20961 18555 20995
rect 22937 20961 22971 20995
rect 23673 20961 23707 20995
rect 27261 20961 27295 20995
rect 32689 20961 32723 20995
rect 34161 20961 34195 20995
rect 36461 20961 36495 20995
rect 38117 20961 38151 20995
rect 1593 20893 1627 20927
rect 5089 20893 5123 20927
rect 5365 20893 5399 20927
rect 6009 20893 6043 20927
rect 6101 20893 6135 20927
rect 6837 20893 6871 20927
rect 7113 20893 7147 20927
rect 8953 20893 8987 20927
rect 9229 20893 9263 20927
rect 9873 20893 9907 20927
rect 10057 20893 10091 20927
rect 10701 20893 10735 20927
rect 10885 20893 10919 20927
rect 11003 20893 11037 20927
rect 11805 20893 11839 20927
rect 12633 20893 12667 20927
rect 14105 20893 14139 20927
rect 16497 20893 16531 20927
rect 19441 20893 19475 20927
rect 19625 20893 19659 20927
rect 19717 20893 19751 20927
rect 20361 20893 20395 20927
rect 20545 20893 20579 20927
rect 23397 20893 23431 20927
rect 23489 20893 23523 20927
rect 26157 20893 26191 20927
rect 26742 20893 26776 20927
rect 27721 20893 27755 20927
rect 28549 20893 28583 20927
rect 28641 20893 28675 20927
rect 29653 20893 29687 20927
rect 29745 20893 29779 20927
rect 30113 20893 30147 20927
rect 33885 20893 33919 20927
rect 36277 20893 36311 20927
rect 5273 20825 5307 20859
rect 8309 20825 8343 20859
rect 9965 20825 9999 20859
rect 10793 20825 10827 20859
rect 11989 20825 12023 20859
rect 13461 20825 13495 20859
rect 14372 20825 14406 20859
rect 18429 20825 18463 20859
rect 19257 20825 19291 20859
rect 22661 20825 22695 20859
rect 28365 20825 28399 20859
rect 32413 20825 32447 20859
rect 35357 20825 35391 20859
rect 35449 20825 35483 20859
rect 9045 20757 9079 20791
rect 12449 20757 12483 20791
rect 15485 20757 15519 20791
rect 17969 20757 18003 20791
rect 18337 20757 18371 20791
rect 20177 20757 20211 20791
rect 23673 20757 23707 20791
rect 24409 20757 24443 20791
rect 26801 20757 26835 20791
rect 35081 20757 35115 20791
rect 35265 20757 35299 20791
rect 5825 20553 5859 20587
rect 9045 20553 9079 20587
rect 11713 20553 11747 20587
rect 13645 20553 13679 20587
rect 14749 20553 14783 20587
rect 16881 20553 16915 20587
rect 21833 20553 21867 20587
rect 22845 20553 22879 20587
rect 26433 20553 26467 20587
rect 27813 20553 27847 20587
rect 28825 20553 28859 20587
rect 33425 20553 33459 20587
rect 6745 20485 6779 20519
rect 6863 20485 6897 20519
rect 8677 20485 8711 20519
rect 8861 20485 8895 20519
rect 9505 20485 9539 20519
rect 12909 20485 12943 20519
rect 14243 20485 14277 20519
rect 14473 20485 14507 20519
rect 15361 20485 15395 20519
rect 15577 20485 15611 20519
rect 16681 20485 16715 20519
rect 29101 20485 29135 20519
rect 37289 20485 37323 20519
rect 2053 20417 2087 20451
rect 4445 20417 4479 20451
rect 4712 20417 4746 20451
rect 6377 20417 6411 20451
rect 6561 20417 6595 20451
rect 6653 20417 6687 20451
rect 7849 20417 7883 20451
rect 7941 20417 7975 20451
rect 9689 20417 9723 20451
rect 10241 20417 10275 20451
rect 10425 20417 10459 20451
rect 11989 20417 12023 20451
rect 13461 20417 13495 20451
rect 14105 20417 14139 20451
rect 14381 20417 14415 20451
rect 14565 20417 14599 20451
rect 17969 20417 18003 20451
rect 18225 20417 18259 20451
rect 20177 20417 20211 20451
rect 21281 20417 21315 20451
rect 22017 20417 22051 20451
rect 22201 20417 22235 20451
rect 22293 20417 22327 20451
rect 22753 20417 22787 20451
rect 26065 20417 26099 20451
rect 27617 20417 27651 20451
rect 27997 20417 28031 20451
rect 28733 20417 28767 20451
rect 28917 20417 28951 20451
rect 30849 20417 30883 20451
rect 31493 20417 31527 20451
rect 33609 20417 33643 20451
rect 33701 20417 33735 20451
rect 34345 20417 34379 20451
rect 34529 20417 34563 20451
rect 36737 20417 36771 20451
rect 37473 20417 37507 20451
rect 37565 20417 37599 20451
rect 7021 20349 7055 20383
rect 8125 20349 8159 20383
rect 11713 20349 11747 20383
rect 11897 20349 11931 20383
rect 19993 20349 20027 20383
rect 20085 20349 20119 20383
rect 20269 20349 20303 20383
rect 23397 20349 23431 20383
rect 23673 20349 23707 20383
rect 25973 20349 26007 20383
rect 26157 20349 26191 20383
rect 26249 20349 26283 20383
rect 27721 20349 27755 20383
rect 28089 20349 28123 20383
rect 28549 20349 28583 20383
rect 30573 20349 30607 20383
rect 32137 20349 32171 20383
rect 33793 20349 33827 20383
rect 36461 20349 36495 20383
rect 12725 20281 12759 20315
rect 15209 20281 15243 20315
rect 25145 20281 25179 20315
rect 31309 20281 31343 20315
rect 34989 20281 35023 20315
rect 37289 20281 37323 20315
rect 1961 20213 1995 20247
rect 7481 20213 7515 20247
rect 10425 20213 10459 20247
rect 15393 20213 15427 20247
rect 16865 20213 16899 20247
rect 17049 20213 17083 20247
rect 19349 20213 19383 20247
rect 19809 20213 19843 20247
rect 21097 20213 21131 20247
rect 27445 20213 27479 20247
rect 32367 20213 32401 20247
rect 34437 20213 34471 20247
rect 6561 20009 6595 20043
rect 12173 20009 12207 20043
rect 15209 20009 15243 20043
rect 16037 20009 16071 20043
rect 16221 20009 16255 20043
rect 16773 20009 16807 20043
rect 18521 20009 18555 20043
rect 19441 20009 19475 20043
rect 23121 20009 23155 20043
rect 27261 20009 27295 20043
rect 27445 20009 27479 20043
rect 31309 20009 31343 20043
rect 32689 20009 32723 20043
rect 35725 20009 35759 20043
rect 19625 19941 19659 19975
rect 23397 19941 23431 19975
rect 33149 19941 33183 19975
rect 1409 19873 1443 19907
rect 1593 19873 1627 19907
rect 1869 19873 1903 19907
rect 7113 19873 7147 19907
rect 7389 19873 7423 19907
rect 13553 19873 13587 19907
rect 14289 19873 14323 19907
rect 14565 19873 14599 19907
rect 15945 19873 15979 19907
rect 18521 19873 18555 19907
rect 20729 19873 20763 19907
rect 31125 19873 31159 19907
rect 37105 19873 37139 19907
rect 37933 19873 37967 19907
rect 38117 19873 38151 19907
rect 6469 19805 6503 19839
rect 6653 19805 6687 19839
rect 8953 19805 8987 19839
rect 10977 19805 11011 19839
rect 11253 19805 11287 19839
rect 13185 19805 13219 19839
rect 13277 19805 13311 19839
rect 14381 19805 14415 19839
rect 14473 19805 14507 19839
rect 15301 19805 15335 19839
rect 15761 19805 15795 19839
rect 16037 19805 16071 19839
rect 16681 19805 16715 19839
rect 16865 19805 16899 19839
rect 17233 19805 17267 19839
rect 17509 19805 17543 19839
rect 18429 19805 18463 19839
rect 18705 19805 18739 19839
rect 22385 19805 22419 19839
rect 23305 19805 23339 19839
rect 23489 19805 23523 19839
rect 23581 19805 23615 19839
rect 24593 19805 24627 19839
rect 25605 19805 25639 19839
rect 25881 19805 25915 19839
rect 28641 19805 28675 19839
rect 28825 19805 28859 19839
rect 29009 19805 29043 19839
rect 29561 19805 29595 19839
rect 29745 19805 29779 19839
rect 30021 19805 30055 19839
rect 30665 19805 30699 19839
rect 31033 19805 31067 19839
rect 32045 19805 32079 19839
rect 32229 19805 32263 19839
rect 32321 19805 32355 19839
rect 32413 19805 32447 19839
rect 33425 19805 33459 19839
rect 35081 19805 35115 19839
rect 35265 19805 35299 19839
rect 35357 19805 35391 19839
rect 35449 19805 35483 19839
rect 9198 19737 9232 19771
rect 12265 19737 12299 19771
rect 19257 19737 19291 19771
rect 19457 19737 19491 19771
rect 27429 19737 27463 19771
rect 27629 19737 27663 19771
rect 10333 19669 10367 19703
rect 10793 19669 10827 19703
rect 11161 19669 11195 19703
rect 13369 19669 13403 19703
rect 13461 19669 13495 19703
rect 14105 19669 14139 19703
rect 18245 19669 18279 19703
rect 24409 19669 24443 19703
rect 29929 19669 29963 19703
rect 30757 19669 30791 19703
rect 30941 19669 30975 19703
rect 33333 19669 33367 19703
rect 33517 19669 33551 19703
rect 33701 19669 33735 19703
rect 7757 19465 7791 19499
rect 9413 19465 9447 19499
rect 9781 19465 9815 19499
rect 9873 19465 9907 19499
rect 10977 19465 11011 19499
rect 13829 19465 13863 19499
rect 14841 19465 14875 19499
rect 16865 19465 16899 19499
rect 18521 19465 18555 19499
rect 18889 19465 18923 19499
rect 26985 19465 27019 19499
rect 27153 19465 27187 19499
rect 32489 19465 32523 19499
rect 34161 19465 34195 19499
rect 36737 19465 36771 19499
rect 12716 19397 12750 19431
rect 15729 19397 15763 19431
rect 15945 19397 15979 19431
rect 19984 19397 20018 19431
rect 22293 19397 22327 19431
rect 26065 19397 26099 19431
rect 27353 19397 27387 19431
rect 31585 19397 31619 19431
rect 32689 19397 32723 19431
rect 34313 19397 34347 19431
rect 34529 19397 34563 19431
rect 37289 19397 37323 19431
rect 6377 19329 6411 19363
rect 6633 19329 6667 19363
rect 8769 19329 8803 19363
rect 10793 19329 10827 19363
rect 11897 19329 11931 19363
rect 14381 19329 14415 19363
rect 14565 19329 14599 19363
rect 14841 19329 14875 19363
rect 15117 19329 15151 19363
rect 16957 19329 16991 19363
rect 17049 19329 17083 19363
rect 17877 19329 17911 19363
rect 18981 19329 19015 19363
rect 23489 19329 23523 19363
rect 25973 19329 26007 19363
rect 26249 19329 26283 19363
rect 28273 19329 28307 19363
rect 28457 19329 28491 19363
rect 28549 19329 28583 19363
rect 29193 19329 29227 19363
rect 30021 19329 30055 19363
rect 31309 19329 31343 19363
rect 33333 19329 33367 19363
rect 34989 19329 35023 19363
rect 37473 19329 37507 19363
rect 37565 19329 37599 19363
rect 1685 19261 1719 19295
rect 1869 19261 1903 19295
rect 2145 19261 2179 19295
rect 10057 19261 10091 19295
rect 12449 19261 12483 19295
rect 16681 19261 16715 19295
rect 19165 19261 19199 19295
rect 19717 19261 19751 19295
rect 22569 19261 22603 19295
rect 23765 19261 23799 19295
rect 28089 19261 28123 19295
rect 29101 19261 29135 19295
rect 29285 19261 29319 19295
rect 29377 19261 29411 19295
rect 30297 19261 30331 19295
rect 31585 19261 31619 19295
rect 33517 19261 33551 19295
rect 35265 19261 35299 19295
rect 8953 19193 8987 19227
rect 11713 19193 11747 19227
rect 17233 19193 17267 19227
rect 37289 19193 37323 19227
rect 15577 19125 15611 19159
rect 15761 19125 15795 19159
rect 18061 19125 18095 19159
rect 21097 19125 21131 19159
rect 25237 19125 25271 19159
rect 25973 19125 26007 19159
rect 27169 19125 27203 19159
rect 29561 19125 29595 19159
rect 31401 19125 31435 19159
rect 32321 19125 32355 19159
rect 32505 19125 32539 19159
rect 33149 19125 33183 19159
rect 34345 19125 34379 19159
rect 1593 18921 1627 18955
rect 2145 18921 2179 18955
rect 6469 18921 6503 18955
rect 10517 18921 10551 18955
rect 10701 18921 10735 18955
rect 16773 18921 16807 18955
rect 19441 18921 19475 18955
rect 21833 18921 21867 18955
rect 22017 18921 22051 18955
rect 26249 18921 26283 18955
rect 27997 18921 28031 18955
rect 28825 18921 28859 18955
rect 29009 18921 29043 18955
rect 30665 18921 30699 18955
rect 31309 18921 31343 18955
rect 34897 18921 34931 18955
rect 35633 18921 35667 18955
rect 14933 18853 14967 18887
rect 23581 18853 23615 18887
rect 9781 18785 9815 18819
rect 10333 18785 10367 18819
rect 11529 18785 11563 18819
rect 11989 18785 12023 18819
rect 16037 18785 16071 18819
rect 17785 18785 17819 18819
rect 17877 18785 17911 18819
rect 26341 18785 26375 18819
rect 27353 18785 27387 18819
rect 37933 18785 37967 18819
rect 2237 18717 2271 18751
rect 6653 18717 6687 18751
rect 8401 18717 8435 18751
rect 9413 18717 9447 18751
rect 9597 18717 9631 18751
rect 10517 18717 10551 18751
rect 11345 18717 11379 18751
rect 12173 18717 12207 18751
rect 12265 18717 12299 18751
rect 13093 18717 13127 18751
rect 13369 18717 13403 18751
rect 15761 18717 15795 18751
rect 17693 18717 17727 18751
rect 17969 18717 18003 18751
rect 19533 18717 19567 18751
rect 21373 18717 21407 18751
rect 22937 18717 22971 18751
rect 23397 18717 23431 18751
rect 25421 18717 25455 18751
rect 25697 18717 25731 18751
rect 26433 18717 26467 18751
rect 27445 18717 27479 18751
rect 30021 18717 30055 18751
rect 30205 18717 30239 18751
rect 30297 18717 30331 18751
rect 30389 18717 30423 18751
rect 32321 18717 32355 18751
rect 32597 18717 32631 18751
rect 33517 18717 33551 18751
rect 34161 18717 34195 18751
rect 35541 18717 35575 18751
rect 10241 18649 10275 18683
rect 14749 18649 14783 18683
rect 16589 18649 16623 18683
rect 16805 18649 16839 18683
rect 21106 18649 21140 18683
rect 21985 18649 22019 18683
rect 22201 18649 22235 18683
rect 24501 18649 24535 18683
rect 26157 18649 26191 18683
rect 28089 18649 28123 18683
rect 28641 18649 28675 18683
rect 28857 18649 28891 18683
rect 31277 18649 31311 18683
rect 31493 18649 31527 18683
rect 33241 18649 33275 18683
rect 33425 18649 33459 18683
rect 34713 18649 34747 18683
rect 37657 18649 37691 18683
rect 8217 18581 8251 18615
rect 11161 18581 11195 18615
rect 11989 18581 12023 18615
rect 12909 18581 12943 18615
rect 13277 18581 13311 18615
rect 15393 18581 15427 18615
rect 15853 18581 15887 18615
rect 16957 18581 16991 18615
rect 18153 18581 18187 18615
rect 19993 18581 20027 18615
rect 22753 18581 22787 18615
rect 24593 18581 24627 18615
rect 25237 18581 25271 18615
rect 25605 18581 25639 18615
rect 26617 18581 26651 18615
rect 31125 18581 31159 18615
rect 32413 18581 32447 18615
rect 32781 18581 32815 18615
rect 33517 18581 33551 18615
rect 33977 18581 34011 18615
rect 34913 18581 34947 18615
rect 35081 18581 35115 18615
rect 36185 18581 36219 18615
rect 10333 18377 10367 18411
rect 10793 18377 10827 18411
rect 12909 18377 12943 18411
rect 16865 18377 16899 18411
rect 19993 18377 20027 18411
rect 21189 18377 21223 18411
rect 24961 18377 24995 18411
rect 25957 18377 25991 18411
rect 29101 18377 29135 18411
rect 31493 18377 31527 18411
rect 33057 18377 33091 18411
rect 33241 18377 33275 18411
rect 37473 18377 37507 18411
rect 10885 18309 10919 18343
rect 26157 18309 26191 18343
rect 26985 18309 27019 18343
rect 31125 18309 31159 18343
rect 31341 18309 31375 18343
rect 8033 18241 8067 18275
rect 8300 18241 8334 18275
rect 10609 18241 10643 18275
rect 11897 18241 11931 18275
rect 13093 18241 13127 18275
rect 14013 18241 14047 18275
rect 15025 18241 15059 18275
rect 19266 18241 19300 18275
rect 19533 18241 19567 18275
rect 20177 18241 20211 18275
rect 20361 18241 20395 18275
rect 21281 18241 21315 18275
rect 21833 18241 21867 18275
rect 24317 18241 24351 18275
rect 25145 18241 25179 18275
rect 25329 18241 25363 18275
rect 27261 18241 27295 18275
rect 28273 18241 28307 18275
rect 29009 18241 29043 18275
rect 29837 18241 29871 18275
rect 32873 18241 32907 18275
rect 32965 18241 32999 18275
rect 36461 18241 36495 18275
rect 37289 18241 37323 18275
rect 37933 18241 37967 18275
rect 10517 18173 10551 18207
rect 10977 18173 11011 18207
rect 11713 18173 11747 18207
rect 11805 18173 11839 18207
rect 11989 18173 12023 18207
rect 13277 18173 13311 18207
rect 14749 18173 14783 18207
rect 22109 18173 22143 18207
rect 26985 18173 27019 18207
rect 30113 18173 30147 18207
rect 34253 18173 34287 18207
rect 34529 18173 34563 18207
rect 9413 18105 9447 18139
rect 14197 18105 14231 18139
rect 17233 18105 17267 18139
rect 23581 18105 23615 18139
rect 32689 18105 32723 18139
rect 1685 18037 1719 18071
rect 11529 18037 11563 18071
rect 16681 18037 16715 18071
rect 16865 18037 16899 18071
rect 18153 18037 18187 18071
rect 24133 18037 24167 18071
rect 25789 18037 25823 18071
rect 25973 18037 26007 18071
rect 27169 18037 27203 18071
rect 28365 18037 28399 18071
rect 31309 18037 31343 18071
rect 36001 18037 36035 18071
rect 36645 18037 36679 18071
rect 38025 18037 38059 18071
rect 14105 17833 14139 17867
rect 16129 17833 16163 17867
rect 18613 17833 18647 17867
rect 19257 17833 19291 17867
rect 19625 17833 19659 17867
rect 23213 17833 23247 17867
rect 24409 17833 24443 17867
rect 25881 17833 25915 17867
rect 26341 17833 26375 17867
rect 30113 17833 30147 17867
rect 32505 17833 32539 17867
rect 34713 17833 34747 17867
rect 35541 17833 35575 17867
rect 13093 17765 13127 17799
rect 21833 17765 21867 17799
rect 25329 17765 25363 17799
rect 32689 17765 32723 17799
rect 33241 17765 33275 17799
rect 35633 17765 35667 17799
rect 1409 17697 1443 17731
rect 2789 17697 2823 17731
rect 9597 17697 9631 17731
rect 10517 17697 10551 17731
rect 14749 17697 14783 17731
rect 17141 17697 17175 17731
rect 18429 17697 18463 17731
rect 19717 17697 19751 17731
rect 26525 17697 26559 17731
rect 37105 17697 37139 17731
rect 37933 17697 37967 17731
rect 38117 17697 38151 17731
rect 8401 17629 8435 17663
rect 9321 17629 9355 17663
rect 10425 17629 10459 17663
rect 10609 17629 10643 17663
rect 10701 17629 10735 17663
rect 11253 17629 11287 17663
rect 11529 17629 11563 17663
rect 12909 17629 12943 17663
rect 14105 17629 14139 17663
rect 14289 17629 14323 17663
rect 17417 17629 17451 17663
rect 18705 17629 18739 17663
rect 19441 17629 19475 17663
rect 20637 17629 20671 17663
rect 21281 17629 21315 17663
rect 21741 17629 21775 17663
rect 22569 17629 22603 17663
rect 23029 17629 23063 17663
rect 23213 17629 23247 17663
rect 23857 17629 23891 17663
rect 24593 17629 24627 17663
rect 26617 17629 26651 17663
rect 26985 17629 27019 17663
rect 27905 17629 27939 17663
rect 28181 17629 28215 17663
rect 28457 17629 28491 17663
rect 28641 17629 28675 17663
rect 31125 17629 31159 17663
rect 33149 17629 33183 17663
rect 33425 17629 33459 17663
rect 34989 17629 35023 17663
rect 35449 17629 35483 17663
rect 35725 17629 35759 17663
rect 1593 17561 1627 17595
rect 9413 17561 9447 17595
rect 12541 17561 12575 17595
rect 12817 17561 12851 17595
rect 15016 17561 15050 17595
rect 18429 17561 18463 17595
rect 22477 17561 22511 17595
rect 25605 17561 25639 17595
rect 30021 17561 30055 17595
rect 32321 17561 32355 17595
rect 33609 17561 33643 17595
rect 34713 17561 34747 17595
rect 8217 17493 8251 17527
rect 8953 17493 8987 17527
rect 10241 17493 10275 17527
rect 12725 17493 12759 17527
rect 20545 17493 20579 17527
rect 21189 17493 21223 17527
rect 23765 17493 23799 17527
rect 25513 17493 25547 17527
rect 25697 17493 25731 17527
rect 26709 17493 26743 17527
rect 26893 17493 26927 17527
rect 27997 17493 28031 17527
rect 31217 17493 31251 17527
rect 32521 17493 32555 17527
rect 34897 17493 34931 17527
rect 1961 17289 1995 17323
rect 9137 17289 9171 17323
rect 10701 17289 10735 17323
rect 10793 17289 10827 17323
rect 14565 17289 14599 17323
rect 15209 17289 15243 17323
rect 16681 17289 16715 17323
rect 18705 17289 18739 17323
rect 22477 17289 22511 17323
rect 27537 17289 27571 17323
rect 32857 17289 32891 17323
rect 33717 17289 33751 17323
rect 33885 17289 33919 17323
rect 37381 17289 37415 17323
rect 13645 17221 13679 17255
rect 16037 17221 16071 17255
rect 27077 17221 27111 17255
rect 33057 17221 33091 17255
rect 33517 17221 33551 17255
rect 35081 17221 35115 17255
rect 38025 17221 38059 17255
rect 2053 17153 2087 17187
rect 7757 17153 7791 17187
rect 8024 17153 8058 17187
rect 9781 17153 9815 17187
rect 10885 17153 10919 17187
rect 11805 17153 11839 17187
rect 13001 17153 13035 17187
rect 13921 17153 13955 17187
rect 14565 17153 14599 17187
rect 14749 17153 14783 17187
rect 15393 17153 15427 17187
rect 15945 17153 15979 17187
rect 16129 17153 16163 17187
rect 17794 17153 17828 17187
rect 18061 17153 18095 17187
rect 18521 17153 18555 17187
rect 18705 17153 18739 17187
rect 22385 17153 22419 17187
rect 24869 17153 24903 17187
rect 25513 17153 25547 17187
rect 25605 17153 25639 17187
rect 25697 17153 25731 17187
rect 25881 17153 25915 17187
rect 27353 17153 27387 17187
rect 28273 17153 28307 17187
rect 37289 17153 37323 17187
rect 37933 17153 37967 17187
rect 9965 17085 9999 17119
rect 10517 17085 10551 17119
rect 11529 17085 11563 17119
rect 13185 17085 13219 17119
rect 13737 17085 13771 17119
rect 19533 17085 19567 17119
rect 19809 17085 19843 17119
rect 24593 17085 24627 17119
rect 27261 17085 27295 17119
rect 27997 17085 28031 17119
rect 31125 17085 31159 17119
rect 31401 17085 31435 17119
rect 34897 17085 34931 17119
rect 36737 17085 36771 17119
rect 10793 17017 10827 17051
rect 14105 17017 14139 17051
rect 25329 17017 25363 17051
rect 29653 17017 29687 17051
rect 9597 16949 9631 16983
rect 12817 16949 12851 16983
rect 13737 16949 13771 16983
rect 21281 16949 21315 16983
rect 23121 16949 23155 16983
rect 27077 16949 27111 16983
rect 32689 16949 32723 16983
rect 32873 16949 32907 16983
rect 33701 16949 33735 16983
rect 10333 16745 10367 16779
rect 16957 16745 16991 16779
rect 24869 16745 24903 16779
rect 26893 16745 26927 16779
rect 31217 16745 31251 16779
rect 32137 16745 32171 16779
rect 33885 16745 33919 16779
rect 34713 16745 34747 16779
rect 35173 16745 35207 16779
rect 22385 16677 22419 16711
rect 23857 16677 23891 16711
rect 27721 16677 27755 16711
rect 31953 16677 31987 16711
rect 34069 16677 34103 16711
rect 8953 16609 8987 16643
rect 11621 16609 11655 16643
rect 11713 16609 11747 16643
rect 12909 16609 12943 16643
rect 13001 16609 13035 16643
rect 15945 16609 15979 16643
rect 19993 16609 20027 16643
rect 20269 16609 20303 16643
rect 22569 16609 22603 16643
rect 25513 16609 25547 16643
rect 26985 16609 27019 16643
rect 28365 16609 28399 16643
rect 28457 16609 28491 16643
rect 28641 16609 28675 16643
rect 30573 16609 30607 16643
rect 34989 16609 35023 16643
rect 36277 16609 36311 16643
rect 11529 16541 11563 16575
rect 13093 16541 13127 16575
rect 14289 16541 14323 16575
rect 14657 16541 14691 16575
rect 15853 16541 15887 16575
rect 16037 16541 16071 16575
rect 16497 16541 16531 16575
rect 16589 16541 16623 16575
rect 16773 16541 16807 16575
rect 17417 16541 17451 16575
rect 18061 16541 18095 16575
rect 19533 16541 19567 16575
rect 22293 16541 22327 16575
rect 23213 16541 23247 16575
rect 23397 16541 23431 16575
rect 23489 16541 23523 16575
rect 23598 16541 23632 16575
rect 24593 16541 24627 16575
rect 24777 16541 24811 16575
rect 24869 16541 24903 16575
rect 25605 16541 25639 16575
rect 26709 16541 26743 16575
rect 26801 16541 26835 16575
rect 27537 16541 27571 16575
rect 28550 16541 28584 16575
rect 30113 16541 30147 16575
rect 30481 16541 30515 16575
rect 31217 16541 31251 16575
rect 31493 16541 31527 16575
rect 32781 16541 32815 16575
rect 33057 16541 33091 16575
rect 34897 16541 34931 16575
rect 35633 16541 35667 16575
rect 9220 16473 9254 16507
rect 14381 16473 14415 16507
rect 14473 16473 14507 16507
rect 22569 16473 22603 16507
rect 31309 16473 31343 16507
rect 32321 16473 32355 16507
rect 32873 16473 32907 16507
rect 33701 16473 33735 16507
rect 35173 16473 35207 16507
rect 36461 16473 36495 16507
rect 38117 16473 38151 16507
rect 11161 16405 11195 16439
rect 13461 16405 13495 16439
rect 14105 16405 14139 16439
rect 17509 16405 17543 16439
rect 18153 16405 18187 16439
rect 19349 16405 19383 16439
rect 21741 16405 21775 16439
rect 25329 16405 25363 16439
rect 25973 16405 26007 16439
rect 28181 16405 28215 16439
rect 30205 16405 30239 16439
rect 30297 16405 30331 16439
rect 30757 16405 30791 16439
rect 32121 16405 32155 16439
rect 33241 16405 33275 16439
rect 33901 16405 33935 16439
rect 35725 16405 35759 16439
rect 9229 16201 9263 16235
rect 12909 16201 12943 16235
rect 15025 16201 15059 16235
rect 20177 16201 20211 16235
rect 23305 16201 23339 16235
rect 29653 16201 29687 16235
rect 30113 16201 30147 16235
rect 32781 16201 32815 16235
rect 37289 16201 37323 16235
rect 38025 16201 38059 16235
rect 10701 16133 10735 16167
rect 10885 16133 10919 16167
rect 23857 16133 23891 16167
rect 32689 16133 32723 16167
rect 34161 16133 34195 16167
rect 36277 16133 36311 16167
rect 9413 16065 9447 16099
rect 11785 16065 11819 16099
rect 13645 16065 13679 16099
rect 13912 16065 13946 16099
rect 15761 16065 15795 16099
rect 17141 16065 17175 16099
rect 20361 16065 20395 16099
rect 21097 16065 21131 16099
rect 22201 16065 22235 16099
rect 22385 16065 22419 16099
rect 23121 16065 23155 16099
rect 24225 16065 24259 16099
rect 24961 16065 24995 16099
rect 25789 16065 25823 16099
rect 26065 16065 26099 16099
rect 27169 16065 27203 16099
rect 27353 16065 27387 16099
rect 27445 16065 27479 16099
rect 27905 16065 27939 16099
rect 30481 16065 30515 16099
rect 31401 16065 31435 16099
rect 34069 16065 34103 16099
rect 34345 16065 34379 16099
rect 37473 16065 37507 16099
rect 37933 16065 37967 16099
rect 11529 15997 11563 16031
rect 17969 15997 18003 16031
rect 18245 15997 18279 16031
rect 22845 15997 22879 16031
rect 25973 15997 26007 16031
rect 30297 15997 30331 16031
rect 30389 15997 30423 16031
rect 33057 15997 33091 16031
rect 36553 15997 36587 16031
rect 25053 15929 25087 15963
rect 34805 15929 34839 15963
rect 2145 15861 2179 15895
rect 15853 15861 15887 15895
rect 17233 15861 17267 15895
rect 19717 15861 19751 15895
rect 21281 15861 21315 15895
rect 22109 15861 22143 15895
rect 22937 15861 22971 15895
rect 25605 15861 25639 15895
rect 27169 15861 27203 15895
rect 28168 15861 28202 15895
rect 31493 15861 31527 15895
rect 32965 15861 32999 15895
rect 33149 15861 33183 15895
rect 34345 15861 34379 15895
rect 10977 15657 11011 15691
rect 13553 15657 13587 15691
rect 18429 15657 18463 15691
rect 20637 15657 20671 15691
rect 24685 15657 24719 15691
rect 28457 15657 28491 15691
rect 29653 15657 29687 15691
rect 35357 15657 35391 15691
rect 11529 15589 11563 15623
rect 14381 15589 14415 15623
rect 19257 15589 19291 15623
rect 22753 15589 22787 15623
rect 26985 15589 27019 15623
rect 1409 15521 1443 15555
rect 3249 15521 3283 15555
rect 14841 15521 14875 15555
rect 16589 15521 16623 15555
rect 19809 15521 19843 15555
rect 20821 15521 20855 15555
rect 25237 15521 25271 15555
rect 25513 15521 25547 15555
rect 27997 15521 28031 15555
rect 30205 15521 30239 15555
rect 31585 15521 31619 15555
rect 32413 15521 32447 15555
rect 32689 15521 32723 15555
rect 35265 15521 35299 15555
rect 37105 15521 37139 15555
rect 10793 15453 10827 15487
rect 11437 15453 11471 15487
rect 11621 15453 11655 15487
rect 12173 15453 12207 15487
rect 17693 15453 17727 15487
rect 17877 15453 17911 15487
rect 18613 15453 18647 15487
rect 20637 15453 20671 15487
rect 20913 15453 20947 15487
rect 22569 15453 22603 15487
rect 23857 15453 23891 15487
rect 24593 15453 24627 15487
rect 28089 15453 28123 15487
rect 28273 15453 28307 15487
rect 29561 15453 29595 15487
rect 29745 15453 29779 15487
rect 30389 15453 30423 15487
rect 30481 15453 30515 15487
rect 30757 15453 30791 15487
rect 31401 15453 31435 15487
rect 35449 15453 35483 15487
rect 35541 15453 35575 15487
rect 38117 15453 38151 15487
rect 3065 15385 3099 15419
rect 12440 15385 12474 15419
rect 14197 15385 14231 15419
rect 15117 15385 15151 15419
rect 21557 15385 21591 15419
rect 21741 15385 21775 15419
rect 23765 15385 23799 15419
rect 37933 15385 37967 15419
rect 17509 15317 17543 15351
rect 19625 15317 19659 15351
rect 19717 15317 19751 15351
rect 20453 15317 20487 15351
rect 21373 15317 21407 15351
rect 30573 15317 30607 15351
rect 31217 15317 31251 15351
rect 34161 15317 34195 15351
rect 2697 15113 2731 15147
rect 13829 15113 13863 15147
rect 15117 15113 15151 15147
rect 19089 15113 19123 15147
rect 20637 15113 20671 15147
rect 23305 15113 23339 15147
rect 24317 15113 24351 15147
rect 25605 15113 25639 15147
rect 26249 15113 26283 15147
rect 29377 15113 29411 15147
rect 29837 15113 29871 15147
rect 30849 15113 30883 15147
rect 32137 15113 32171 15147
rect 32305 15113 32339 15147
rect 12633 15045 12667 15079
rect 13369 15045 13403 15079
rect 18889 15045 18923 15079
rect 20913 15045 20947 15079
rect 24133 15045 24167 15079
rect 25697 15045 25731 15079
rect 31012 15045 31046 15079
rect 31217 15045 31251 15079
rect 32505 15045 32539 15079
rect 33333 15045 33367 15079
rect 35541 15045 35575 15079
rect 36645 15045 36679 15079
rect 2789 14977 2823 15011
rect 3433 14977 3467 15011
rect 12817 14977 12851 15011
rect 14381 14977 14415 15011
rect 15209 14977 15243 15011
rect 15669 14977 15703 15011
rect 19717 14977 19751 15011
rect 19901 14977 19935 15011
rect 20821 14977 20855 15011
rect 21005 14977 21039 15011
rect 21123 14977 21157 15011
rect 23121 14977 23155 15011
rect 23305 14977 23339 15011
rect 24409 14977 24443 15011
rect 24869 14977 24903 15011
rect 25053 14977 25087 15011
rect 26249 14977 26283 15011
rect 26433 14977 26467 15011
rect 27721 14977 27755 15011
rect 29193 14977 29227 15011
rect 30021 14977 30055 15011
rect 30297 14977 30331 15011
rect 33057 14977 33091 15011
rect 35449 14977 35483 15011
rect 35725 14977 35759 15011
rect 36553 14977 36587 15011
rect 37473 14977 37507 15011
rect 16681 14909 16715 14943
rect 16957 14909 16991 14943
rect 18429 14909 18463 14943
rect 21281 14909 21315 14943
rect 21833 14909 21867 14943
rect 22109 14909 22143 14943
rect 24961 14909 24995 14943
rect 27537 14909 27571 14943
rect 27629 14909 27663 14943
rect 29009 14909 29043 14943
rect 30205 14909 30239 14943
rect 34805 14909 34839 14943
rect 13645 14841 13679 14875
rect 15853 14841 15887 14875
rect 19257 14841 19291 14875
rect 1869 14773 1903 14807
rect 3341 14773 3375 14807
rect 14473 14773 14507 14807
rect 19073 14773 19107 14807
rect 19717 14773 19751 14807
rect 24133 14773 24167 14807
rect 28089 14773 28123 14807
rect 30297 14773 30331 14807
rect 31033 14773 31067 14807
rect 32321 14773 32355 14807
rect 35725 14773 35759 14807
rect 37565 14773 37599 14807
rect 13001 14569 13035 14603
rect 17325 14569 17359 14603
rect 17693 14569 17727 14603
rect 21649 14569 21683 14603
rect 31677 14569 31711 14603
rect 33793 14569 33827 14603
rect 16865 14501 16899 14535
rect 21097 14501 21131 14535
rect 24409 14501 24443 14535
rect 35357 14501 35391 14535
rect 3065 14433 3099 14467
rect 20545 14433 20579 14467
rect 22569 14433 22603 14467
rect 23581 14433 23615 14467
rect 26157 14433 26191 14467
rect 27077 14433 27111 14467
rect 28825 14433 28859 14467
rect 29561 14433 29595 14467
rect 29837 14433 29871 14467
rect 31125 14433 31159 14467
rect 32413 14433 32447 14467
rect 36461 14433 36495 14467
rect 38117 14433 38151 14467
rect 1409 14365 1443 14399
rect 3249 14365 3283 14399
rect 3801 14365 3835 14399
rect 13185 14365 13219 14399
rect 14749 14365 14783 14399
rect 15761 14365 15795 14399
rect 15945 14365 15979 14399
rect 16589 14365 16623 14399
rect 17509 14365 17543 14399
rect 17785 14365 17819 14399
rect 18245 14365 18279 14399
rect 18429 14365 18463 14399
rect 19625 14365 19659 14399
rect 20453 14365 20487 14399
rect 20637 14365 20671 14399
rect 21281 14365 21315 14399
rect 22201 14365 22235 14399
rect 22477 14365 22511 14399
rect 23397 14365 23431 14399
rect 31309 14365 31343 14399
rect 32137 14365 32171 14399
rect 36277 14365 36311 14399
rect 33747 14331 33781 14365
rect 16865 14297 16899 14331
rect 22109 14297 22143 14331
rect 25881 14297 25915 14331
rect 27353 14297 27387 14331
rect 31493 14297 31527 14331
rect 33977 14297 34011 14331
rect 35173 14297 35207 14331
rect 14657 14229 14691 14263
rect 15945 14229 15979 14263
rect 16681 14229 16715 14263
rect 18337 14229 18371 14263
rect 19533 14229 19567 14263
rect 21373 14229 21407 14263
rect 21465 14229 21499 14263
rect 22753 14229 22787 14263
rect 23213 14229 23247 14263
rect 31401 14229 31435 14263
rect 33609 14229 33643 14263
rect 12633 14025 12667 14059
rect 17601 14025 17635 14059
rect 22201 14025 22235 14059
rect 25329 14025 25363 14059
rect 27813 14025 27847 14059
rect 28457 14025 28491 14059
rect 31033 14025 31067 14059
rect 31401 14025 31435 14059
rect 34989 14025 35023 14059
rect 37565 14025 37599 14059
rect 13369 13957 13403 13991
rect 17233 13957 17267 13991
rect 17417 13957 17451 13991
rect 21833 13957 21867 13991
rect 27445 13957 27479 13991
rect 27661 13957 27695 13991
rect 22063 13923 22097 13957
rect 1869 13889 1903 13923
rect 12725 13889 12759 13923
rect 13921 13889 13955 13923
rect 18429 13889 18463 13923
rect 18521 13889 18555 13923
rect 18705 13889 18739 13923
rect 19901 13889 19935 13923
rect 20637 13889 20671 13923
rect 20729 13889 20763 13923
rect 20913 13889 20947 13923
rect 22937 13889 22971 13923
rect 25513 13889 25547 13923
rect 26157 13889 26191 13923
rect 30205 13889 30239 13923
rect 31217 13889 31251 13923
rect 31309 13889 31343 13923
rect 32505 13889 32539 13923
rect 32781 13889 32815 13923
rect 33793 13889 33827 13923
rect 34069 13889 34103 13923
rect 34161 13889 34195 13923
rect 36737 13889 36771 13923
rect 37473 13889 37507 13923
rect 2053 13821 2087 13855
rect 2789 13821 2823 13855
rect 13185 13821 13219 13855
rect 14197 13821 14231 13855
rect 15669 13821 15703 13855
rect 18245 13821 18279 13855
rect 18613 13821 18647 13855
rect 23213 13821 23247 13855
rect 24685 13821 24719 13855
rect 29929 13821 29963 13855
rect 31585 13821 31619 13855
rect 33885 13821 33919 13855
rect 34345 13821 34379 13855
rect 36461 13821 36495 13855
rect 19717 13753 19751 13787
rect 20453 13685 20487 13719
rect 20637 13685 20671 13719
rect 22017 13685 22051 13719
rect 26341 13685 26375 13719
rect 27629 13685 27663 13719
rect 2513 13481 2547 13515
rect 16865 13481 16899 13515
rect 18061 13481 18095 13515
rect 20361 13481 20395 13515
rect 21741 13481 21775 13515
rect 23213 13481 23247 13515
rect 24961 13481 24995 13515
rect 27813 13481 27847 13515
rect 29653 13481 29687 13515
rect 30021 13481 30055 13515
rect 33701 13481 33735 13515
rect 34161 13481 34195 13515
rect 21925 13413 21959 13447
rect 34713 13413 34747 13447
rect 16405 13345 16439 13379
rect 17325 13345 17359 13379
rect 17509 13345 17543 13379
rect 21005 13345 21039 13379
rect 29561 13345 29595 13379
rect 30941 13345 30975 13379
rect 31309 13345 31343 13379
rect 32873 13345 32907 13379
rect 35081 13345 35115 13379
rect 38117 13345 38151 13379
rect 1593 13277 1627 13311
rect 2605 13277 2639 13311
rect 17233 13277 17267 13311
rect 18613 13277 18647 13311
rect 19625 13277 19659 13311
rect 20821 13277 20855 13311
rect 22477 13277 22511 13311
rect 22661 13277 22695 13311
rect 23397 13277 23431 13311
rect 24869 13277 24903 13311
rect 26249 13277 26283 13311
rect 26433 13277 26467 13311
rect 26893 13277 26927 13311
rect 27629 13277 27663 13311
rect 29837 13277 29871 13311
rect 31125 13277 31159 13311
rect 32597 13277 32631 13311
rect 33885 13277 33919 13311
rect 33977 13277 34011 13311
rect 34161 13277 34195 13311
rect 34897 13277 34931 13311
rect 35541 13277 35575 13311
rect 36277 13277 36311 13311
rect 16129 13209 16163 13243
rect 18245 13209 18279 13243
rect 18429 13209 18463 13243
rect 21557 13209 21591 13243
rect 21773 13209 21807 13243
rect 25605 13209 25639 13243
rect 28825 13209 28859 13243
rect 29009 13209 29043 13243
rect 35633 13209 35667 13243
rect 35817 13209 35851 13243
rect 36461 13209 36495 13243
rect 14657 13141 14691 13175
rect 18337 13141 18371 13175
rect 19809 13141 19843 13175
rect 20729 13141 20763 13175
rect 22661 13141 22695 13175
rect 25697 13141 25731 13175
rect 26341 13141 26375 13175
rect 27077 13141 27111 13175
rect 35718 13141 35752 13175
rect 15393 12937 15427 12971
rect 18797 12937 18831 12971
rect 24869 12937 24903 12971
rect 31493 12937 31527 12971
rect 32295 12937 32329 12971
rect 34411 12937 34445 12971
rect 35909 12937 35943 12971
rect 37657 12937 37691 12971
rect 14657 12869 14691 12903
rect 14841 12869 14875 12903
rect 19073 12869 19107 12903
rect 19165 12869 19199 12903
rect 21005 12869 21039 12903
rect 21189 12869 21223 12903
rect 22385 12869 22419 12903
rect 24777 12869 24811 12903
rect 26985 12869 27019 12903
rect 27169 12869 27203 12903
rect 28641 12869 28675 12903
rect 28825 12869 28859 12903
rect 32505 12869 32539 12903
rect 34621 12869 34655 12903
rect 36553 12869 36587 12903
rect 2053 12801 2087 12835
rect 14105 12801 14139 12835
rect 15577 12801 15611 12835
rect 16957 12801 16991 12835
rect 18981 12801 19015 12835
rect 19303 12801 19337 12835
rect 19439 12823 19473 12857
rect 20085 12801 20119 12835
rect 22109 12801 22143 12835
rect 22293 12801 22327 12835
rect 22569 12801 22603 12835
rect 22845 12801 22879 12835
rect 23397 12801 23431 12835
rect 24225 12801 24259 12835
rect 25605 12801 25639 12835
rect 26249 12801 26283 12835
rect 26433 12801 26467 12835
rect 27905 12801 27939 12835
rect 29561 12801 29595 12835
rect 29745 12801 29779 12835
rect 29929 12801 29963 12835
rect 31033 12801 31067 12835
rect 31217 12801 31251 12835
rect 35357 12801 35391 12835
rect 35817 12801 35851 12835
rect 36001 12801 36035 12835
rect 36645 12801 36679 12835
rect 37565 12801 37599 12835
rect 17233 12733 17267 12767
rect 20269 12733 20303 12767
rect 25421 12733 25455 12767
rect 29653 12733 29687 12767
rect 31125 12733 31159 12767
rect 31309 12733 31343 12767
rect 33517 12733 33551 12767
rect 33793 12733 33827 12767
rect 35081 12733 35115 12767
rect 35265 12733 35299 12767
rect 34253 12665 34287 12699
rect 1961 12597 1995 12631
rect 14013 12597 14047 12631
rect 23489 12597 23523 12631
rect 24133 12597 24167 12631
rect 25789 12597 25823 12631
rect 26341 12597 26375 12631
rect 27721 12597 27755 12631
rect 29469 12597 29503 12631
rect 32137 12597 32171 12631
rect 32321 12597 32355 12631
rect 34437 12597 34471 12631
rect 35173 12597 35207 12631
rect 18061 12393 18095 12427
rect 24409 12393 24443 12427
rect 25697 12393 25731 12427
rect 28825 12393 28859 12427
rect 29653 12393 29687 12427
rect 31033 12393 31067 12427
rect 33701 12393 33735 12427
rect 34897 12393 34931 12427
rect 35725 12393 35759 12427
rect 21649 12325 21683 12359
rect 30481 12325 30515 12359
rect 1409 12257 1443 12291
rect 1593 12257 1627 12291
rect 2789 12257 2823 12291
rect 14197 12257 14231 12291
rect 17509 12257 17543 12291
rect 19349 12257 19383 12291
rect 19809 12257 19843 12291
rect 25053 12257 25087 12291
rect 32229 12257 32263 12291
rect 32413 12257 32447 12291
rect 15945 12189 15979 12223
rect 17233 12189 17267 12223
rect 18245 12189 18279 12223
rect 18429 12189 18463 12223
rect 19441 12189 19475 12223
rect 20453 12189 20487 12223
rect 20637 12189 20671 12223
rect 20821 12189 20855 12223
rect 21557 12189 21591 12223
rect 21925 12189 21959 12223
rect 22385 12189 22419 12223
rect 23029 12189 23063 12223
rect 23673 12189 23707 12223
rect 23857 12189 23891 12223
rect 25605 12189 25639 12223
rect 25881 12189 25915 12223
rect 26617 12189 26651 12223
rect 29009 12189 29043 12223
rect 29745 12189 29779 12223
rect 30205 12189 30239 12223
rect 30481 12189 30515 12223
rect 30941 12189 30975 12223
rect 31309 12189 31343 12223
rect 33517 12189 33551 12223
rect 33793 12189 33827 12223
rect 34989 12189 35023 12223
rect 35817 12189 35851 12223
rect 36277 12189 36311 12223
rect 15669 12121 15703 12155
rect 18613 12121 18647 12155
rect 20545 12121 20579 12155
rect 23213 12121 23247 12155
rect 23765 12121 23799 12155
rect 24869 12121 24903 12155
rect 26065 12121 26099 12155
rect 26893 12121 26927 12155
rect 31217 12121 31251 12155
rect 36461 12121 36495 12155
rect 38117 12121 38151 12155
rect 16865 12053 16899 12087
rect 17325 12053 17359 12087
rect 18337 12053 18371 12087
rect 20269 12053 20303 12087
rect 24777 12053 24811 12087
rect 28365 12053 28399 12087
rect 30297 12053 30331 12087
rect 31125 12053 31159 12087
rect 31769 12053 31803 12087
rect 32137 12053 32171 12087
rect 33333 12053 33367 12087
rect 17233 11849 17267 11883
rect 17693 11849 17727 11883
rect 17861 11849 17895 11883
rect 18613 11849 18647 11883
rect 21281 11849 21315 11883
rect 25789 11849 25823 11883
rect 26157 11849 26191 11883
rect 30941 11849 30975 11883
rect 32137 11849 32171 11883
rect 36093 11849 36127 11883
rect 37657 11849 37691 11883
rect 15393 11781 15427 11815
rect 18061 11781 18095 11815
rect 22017 11781 22051 11815
rect 25697 11781 25731 11815
rect 29469 11781 29503 11815
rect 32289 11781 32323 11815
rect 32505 11781 32539 11815
rect 34621 11781 34655 11815
rect 12909 11713 12943 11747
rect 15577 11713 15611 11747
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 18521 11713 18555 11747
rect 18705 11713 18739 11747
rect 19809 11713 19843 11747
rect 20821 11713 20855 11747
rect 21097 11713 21131 11747
rect 21833 11713 21867 11747
rect 31401 11713 31435 11747
rect 32965 11713 32999 11747
rect 36737 11713 36771 11747
rect 37749 11713 37783 11747
rect 1593 11645 1627 11679
rect 1777 11645 1811 11679
rect 2053 11645 2087 11679
rect 13185 11645 13219 11679
rect 20085 11645 20119 11679
rect 21005 11645 21039 11679
rect 22845 11645 22879 11679
rect 23121 11645 23155 11679
rect 25605 11645 25639 11679
rect 26985 11645 27019 11679
rect 27261 11645 27295 11679
rect 29193 11645 29227 11679
rect 34345 11645 34379 11679
rect 14657 11509 14691 11543
rect 17877 11509 17911 11543
rect 20821 11509 20855 11543
rect 22201 11509 22235 11543
rect 24593 11509 24627 11543
rect 28733 11509 28767 11543
rect 31585 11509 31619 11543
rect 32321 11509 32355 11543
rect 33057 11509 33091 11543
rect 33885 11509 33919 11543
rect 36645 11509 36679 11543
rect 1961 11305 1995 11339
rect 14197 11305 14231 11339
rect 14933 11305 14967 11339
rect 17601 11305 17635 11339
rect 19441 11305 19475 11339
rect 22661 11305 22695 11339
rect 26801 11305 26835 11339
rect 27537 11305 27571 11339
rect 29653 11305 29687 11339
rect 30205 11305 30239 11339
rect 34161 11305 34195 11339
rect 35081 11305 35115 11339
rect 19257 11237 19291 11271
rect 35725 11237 35759 11271
rect 16681 11169 16715 11203
rect 18245 11169 18279 11203
rect 18705 11169 18739 11203
rect 21465 11169 21499 11203
rect 22845 11169 22879 11203
rect 24409 11169 24443 11203
rect 24685 11169 24719 11203
rect 25697 11169 25731 11203
rect 26065 11169 26099 11203
rect 28089 11169 28123 11203
rect 31953 11169 31987 11203
rect 32413 11169 32447 11203
rect 32689 11169 32723 11203
rect 36277 11169 36311 11203
rect 2053 11101 2087 11135
rect 14289 11101 14323 11135
rect 17325 11101 17359 11135
rect 18061 11101 18095 11135
rect 18337 11101 18371 11135
rect 19441 11101 19475 11135
rect 19625 11101 19659 11135
rect 20729 11101 20763 11135
rect 21005 11101 21039 11135
rect 21833 11101 21867 11135
rect 21961 11101 21995 11135
rect 22661 11101 22695 11135
rect 22937 11101 22971 11135
rect 23581 11101 23615 11135
rect 25881 11101 25915 11135
rect 25973 11101 26007 11135
rect 26157 11101 26191 11135
rect 26893 11101 26927 11135
rect 27445 11101 27479 11135
rect 28365 11101 28399 11135
rect 29745 11101 29779 11135
rect 34989 11101 35023 11135
rect 35817 11101 35851 11135
rect 16405 11033 16439 11067
rect 17601 11033 17635 11067
rect 21649 11033 21683 11067
rect 21741 11033 21775 11067
rect 31677 11033 31711 11067
rect 36461 11033 36495 11067
rect 38117 11033 38151 11067
rect 17417 10965 17451 10999
rect 22477 10965 22511 10999
rect 23765 10965 23799 10999
rect 14105 10761 14139 10795
rect 14933 10761 14967 10795
rect 17233 10761 17267 10795
rect 17969 10761 18003 10795
rect 18337 10761 18371 10795
rect 19625 10761 19659 10795
rect 21281 10761 21315 10795
rect 22569 10761 22603 10795
rect 24501 10761 24535 10795
rect 27353 10761 27387 10795
rect 29193 10761 29227 10795
rect 30573 10761 30607 10795
rect 33885 10761 33919 10795
rect 17141 10693 17175 10727
rect 17785 10693 17819 10727
rect 18153 10693 18187 10727
rect 22661 10693 22695 10727
rect 24133 10693 24167 10727
rect 24333 10693 24367 10727
rect 25145 10693 25179 10727
rect 25329 10693 25363 10727
rect 26157 10693 26191 10727
rect 31125 10693 31159 10727
rect 31309 10693 31343 10727
rect 36553 10693 36587 10727
rect 1593 10625 1627 10659
rect 14197 10625 14231 10659
rect 14841 10625 14875 10659
rect 15761 10625 15795 10659
rect 15945 10625 15979 10659
rect 18061 10625 18095 10659
rect 18981 10625 19015 10659
rect 19165 10625 19199 10659
rect 19809 10625 19843 10659
rect 20821 10625 20855 10659
rect 21097 10625 21131 10659
rect 22753 10625 22787 10659
rect 23397 10625 23431 10659
rect 23581 10625 23615 10659
rect 25237 10625 25271 10659
rect 27261 10625 27295 10659
rect 28733 10625 28767 10659
rect 29377 10625 29411 10659
rect 29745 10625 29779 10659
rect 30389 10625 30423 10659
rect 32137 10625 32171 10659
rect 37381 10625 37415 10659
rect 15669 10557 15703 10591
rect 15853 10557 15887 10591
rect 21005 10557 21039 10591
rect 23489 10557 23523 10591
rect 28457 10557 28491 10591
rect 29837 10557 29871 10591
rect 32413 10557 32447 10591
rect 35817 10557 35851 10591
rect 36737 10557 36771 10591
rect 19073 10489 19107 10523
rect 22385 10489 22419 10523
rect 24961 10489 24995 10523
rect 25513 10489 25547 10523
rect 15485 10421 15519 10455
rect 20821 10421 20855 10455
rect 22937 10421 22971 10455
rect 24317 10421 24351 10455
rect 26065 10421 26099 10455
rect 29377 10421 29411 10455
rect 37473 10421 37507 10455
rect 17325 10217 17359 10251
rect 18337 10217 18371 10251
rect 19717 10217 19751 10251
rect 19993 10217 20027 10251
rect 20545 10217 20579 10251
rect 21097 10217 21131 10251
rect 22937 10217 22971 10251
rect 23581 10217 23615 10251
rect 27537 10217 27571 10251
rect 27813 10217 27847 10251
rect 30941 10217 30975 10251
rect 31677 10217 31711 10251
rect 32229 10217 32263 10251
rect 34989 10217 35023 10251
rect 35633 10217 35667 10251
rect 22201 10149 22235 10183
rect 17969 10081 18003 10115
rect 20821 10081 20855 10115
rect 22753 10081 22787 10115
rect 24961 10081 24995 10115
rect 28181 10081 28215 10115
rect 34161 10081 34195 10115
rect 36277 10081 36311 10115
rect 36461 10081 36495 10115
rect 38117 10081 38151 10115
rect 14105 10013 14139 10047
rect 14933 10013 14967 10047
rect 16037 10013 16071 10047
rect 16313 10013 16347 10047
rect 16865 10013 16899 10047
rect 16957 10013 16991 10047
rect 17325 10013 17359 10047
rect 18153 10013 18187 10047
rect 19349 10013 19383 10047
rect 19441 10013 19475 10047
rect 19809 10013 19843 10047
rect 20913 10013 20947 10047
rect 23581 10013 23615 10047
rect 23673 10013 23707 10047
rect 23857 10013 23891 10047
rect 27721 10013 27755 10047
rect 28089 10013 28123 10047
rect 28733 10013 28767 10047
rect 28825 10013 28859 10047
rect 29837 10013 29871 10047
rect 30849 10013 30883 10047
rect 31493 10013 31527 10047
rect 32137 10013 32171 10047
rect 34897 10013 34931 10047
rect 35541 10013 35575 10047
rect 20453 9945 20487 9979
rect 22201 9945 22235 9979
rect 25237 9945 25271 9979
rect 29009 9945 29043 9979
rect 14197 9877 14231 9911
rect 14841 9877 14875 9911
rect 17509 9877 17543 9911
rect 22661 9877 22695 9911
rect 23397 9877 23431 9911
rect 26709 9877 26743 9911
rect 28733 9877 28767 9911
rect 29653 9877 29687 9911
rect 18061 9673 18095 9707
rect 18245 9673 18279 9707
rect 19073 9673 19107 9707
rect 20821 9673 20855 9707
rect 22109 9673 22143 9707
rect 25421 9673 25455 9707
rect 30389 9673 30423 9707
rect 17877 9605 17911 9639
rect 18153 9605 18187 9639
rect 21281 9605 21315 9639
rect 22753 9605 22787 9639
rect 27537 9605 27571 9639
rect 27629 9605 27663 9639
rect 27905 9605 27939 9639
rect 28917 9605 28951 9639
rect 30941 9605 30975 9639
rect 36645 9605 36679 9639
rect 13093 9537 13127 9571
rect 15853 9537 15887 9571
rect 16681 9537 16715 9571
rect 17141 9537 17175 9571
rect 18889 9537 18923 9571
rect 18981 9537 19015 9571
rect 19717 9537 19751 9571
rect 20177 9537 20211 9571
rect 21005 9537 21039 9571
rect 23673 9537 23707 9571
rect 24041 9537 24075 9571
rect 24133 9537 24167 9571
rect 25237 9537 25271 9571
rect 26065 9537 26099 9571
rect 27261 9537 27295 9571
rect 27419 9537 27453 9571
rect 27721 9537 27755 9571
rect 31033 9537 31067 9571
rect 35817 9537 35851 9571
rect 36737 9537 36771 9571
rect 37473 9537 37507 9571
rect 13369 9469 13403 9503
rect 16129 9469 16163 9503
rect 16957 9469 16991 9503
rect 19257 9469 19291 9503
rect 19993 9469 20027 9503
rect 21189 9469 21223 9503
rect 22385 9469 22419 9503
rect 24961 9469 24995 9503
rect 25973 9469 26007 9503
rect 26157 9469 26191 9503
rect 26249 9469 26283 9503
rect 28641 9469 28675 9503
rect 35173 9469 35207 9503
rect 18429 9401 18463 9435
rect 19165 9401 19199 9435
rect 20361 9401 20395 9435
rect 26433 9401 26467 9435
rect 34161 9401 34195 9435
rect 1593 9333 1627 9367
rect 2881 9333 2915 9367
rect 14841 9333 14875 9367
rect 16773 9333 16807 9367
rect 17325 9333 17359 9367
rect 19993 9333 20027 9367
rect 21005 9333 21039 9367
rect 22477 9333 22511 9367
rect 22615 9333 22649 9367
rect 23489 9333 23523 9367
rect 23673 9333 23707 9367
rect 25053 9333 25087 9367
rect 37565 9333 37599 9367
rect 13461 9129 13495 9163
rect 14105 9129 14139 9163
rect 16405 9129 16439 9163
rect 17601 9129 17635 9163
rect 21465 9129 21499 9163
rect 21649 9129 21683 9163
rect 22293 9129 22327 9163
rect 22753 9129 22787 9163
rect 23673 9129 23707 9163
rect 29653 9129 29687 9163
rect 31217 9129 31251 9163
rect 35449 9129 35483 9163
rect 18521 9061 18555 9095
rect 19533 9061 19567 9095
rect 24961 9061 24995 9095
rect 30573 9061 30607 9095
rect 1409 8993 1443 9027
rect 1869 8993 1903 9027
rect 15577 8993 15611 9027
rect 15853 8993 15887 9027
rect 17141 8993 17175 9027
rect 21281 8993 21315 9027
rect 25973 8993 26007 9027
rect 26257 8993 26291 9027
rect 37197 8993 37231 9027
rect 37933 8993 37967 9027
rect 3985 8925 4019 8959
rect 4629 8925 4663 8959
rect 13553 8925 13587 8959
rect 16497 8925 16531 8959
rect 17233 8925 17267 8959
rect 17601 8925 17635 8959
rect 18245 8925 18279 8959
rect 19257 8925 19291 8959
rect 20177 8925 20211 8959
rect 21189 8925 21223 8959
rect 21465 8925 21499 8959
rect 22201 8925 22235 8959
rect 22569 8925 22603 8959
rect 23673 8925 23707 8959
rect 23857 8925 23891 8959
rect 26065 8925 26099 8959
rect 26157 8925 26191 8959
rect 27169 8925 27203 8959
rect 27905 8925 27939 8959
rect 28181 8925 28215 8959
rect 29561 8925 29595 8959
rect 29837 8925 29871 8959
rect 30665 8925 30699 8959
rect 31125 8925 31159 8959
rect 38117 8925 38151 8959
rect 1593 8857 1627 8891
rect 18337 8857 18371 8891
rect 18521 8857 18555 8891
rect 19533 8857 19567 8891
rect 24593 8857 24627 8891
rect 24777 8857 24811 8891
rect 26893 8857 26927 8891
rect 27077 8857 27111 8891
rect 27445 8857 27479 8891
rect 30021 8857 30055 8891
rect 3893 8789 3927 8823
rect 17785 8789 17819 8823
rect 19349 8789 19383 8823
rect 20269 8789 20303 8823
rect 24409 8789 24443 8823
rect 24685 8789 24719 8823
rect 26433 8789 26467 8823
rect 27261 8789 27295 8823
rect 1961 8585 1995 8619
rect 14841 8585 14875 8619
rect 16681 8585 16715 8619
rect 17969 8585 18003 8619
rect 18153 8585 18187 8619
rect 20453 8585 20487 8619
rect 22845 8585 22879 8619
rect 23949 8585 23983 8619
rect 24317 8585 24351 8619
rect 24869 8585 24903 8619
rect 4353 8517 4387 8551
rect 17785 8517 17819 8551
rect 18781 8517 18815 8551
rect 18981 8517 19015 8551
rect 19809 8517 19843 8551
rect 21097 8517 21131 8551
rect 23765 8517 23799 8551
rect 24041 8517 24075 8551
rect 25053 8517 25087 8551
rect 29009 8517 29043 8551
rect 2053 8449 2087 8483
rect 5181 8449 5215 8483
rect 15209 8449 15243 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 17141 8449 17175 8483
rect 17877 8449 17911 8483
rect 19625 8449 19659 8483
rect 20361 8449 20395 8483
rect 21281 8449 21315 8483
rect 22017 8449 22051 8483
rect 22753 8449 22787 8483
rect 22937 8449 22971 8483
rect 24133 8449 24167 8483
rect 24777 8449 24811 8483
rect 25145 8449 25179 8483
rect 26157 8449 26191 8483
rect 27445 8449 27479 8483
rect 36737 8449 36771 8483
rect 37841 8449 37875 8483
rect 2881 8381 2915 8415
rect 4537 8381 4571 8415
rect 15301 8381 15335 8415
rect 15485 8381 15519 8415
rect 19441 8381 19475 8415
rect 24961 8381 24995 8415
rect 26433 8381 26467 8415
rect 27721 8381 27755 8415
rect 28733 8381 28767 8415
rect 30481 8381 30515 8415
rect 5089 8313 5123 8347
rect 17601 8313 17635 8347
rect 18613 8245 18647 8279
rect 18797 8245 18831 8279
rect 22201 8245 22235 8279
rect 15485 8041 15519 8075
rect 18429 8041 18463 8075
rect 19625 8041 19659 8075
rect 22201 8041 22235 8075
rect 23673 8041 23707 8075
rect 30297 8041 30331 8075
rect 30941 8041 30975 8075
rect 38117 8041 38151 8075
rect 17417 7973 17451 8007
rect 22937 7973 22971 8007
rect 23857 7973 23891 8007
rect 3985 7905 4019 7939
rect 5641 7905 5675 7939
rect 5825 7905 5859 7939
rect 26157 7905 26191 7939
rect 26249 7905 26283 7939
rect 1777 7837 1811 7871
rect 15393 7837 15427 7871
rect 15577 7837 15611 7871
rect 16221 7837 16255 7871
rect 16405 7837 16439 7871
rect 17049 7837 17083 7871
rect 17233 7837 17267 7871
rect 18245 7837 18279 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 22385 7837 22419 7871
rect 24961 7837 24995 7871
rect 25973 7837 26007 7871
rect 26065 7837 26099 7871
rect 26893 7837 26927 7871
rect 27031 7837 27065 7871
rect 27169 7837 27203 7871
rect 27353 7837 27387 7871
rect 28181 7837 28215 7871
rect 28365 7837 28399 7871
rect 28549 7837 28583 7871
rect 29561 7837 29595 7871
rect 30205 7837 30239 7871
rect 31033 7837 31067 7871
rect 34989 7837 35023 7871
rect 35633 7837 35667 7871
rect 17877 7769 17911 7803
rect 18061 7769 18095 7803
rect 18153 7769 18187 7803
rect 19609 7769 19643 7803
rect 19809 7769 19843 7803
rect 22937 7769 22971 7803
rect 23489 7769 23523 7803
rect 23705 7769 23739 7803
rect 25053 7769 25087 7803
rect 25329 7769 25363 7803
rect 27261 7769 27295 7803
rect 27997 7769 28031 7803
rect 29653 7769 29687 7803
rect 35081 7769 35115 7803
rect 35817 7769 35851 7803
rect 37473 7769 37507 7803
rect 16037 7701 16071 7735
rect 19441 7701 19475 7735
rect 22477 7701 22511 7735
rect 24777 7701 24811 7735
rect 25145 7701 25179 7735
rect 26433 7701 26467 7735
rect 27537 7701 27571 7735
rect 28273 7701 28307 7735
rect 15761 7497 15795 7531
rect 20085 7497 20119 7531
rect 22201 7497 22235 7531
rect 23397 7497 23431 7531
rect 26341 7497 26375 7531
rect 27169 7497 27203 7531
rect 15853 7429 15887 7463
rect 17969 7429 18003 7463
rect 18185 7429 18219 7463
rect 20913 7429 20947 7463
rect 21005 7429 21039 7463
rect 28549 7429 28583 7463
rect 1777 7361 1811 7395
rect 19257 7361 19291 7395
rect 19441 7361 19475 7395
rect 19533 7361 19567 7395
rect 19993 7361 20027 7395
rect 20177 7361 20211 7395
rect 20821 7361 20855 7395
rect 21123 7361 21157 7395
rect 22017 7361 22051 7395
rect 22845 7361 22879 7395
rect 23213 7361 23247 7395
rect 24041 7361 24075 7395
rect 24685 7361 24719 7395
rect 24961 7361 24995 7395
rect 25145 7361 25179 7395
rect 25973 7361 26007 7395
rect 26157 7361 26191 7395
rect 27166 7361 27200 7395
rect 27629 7361 27663 7395
rect 35633 7361 35667 7395
rect 1961 7293 1995 7327
rect 2789 7293 2823 7327
rect 16037 7293 16071 7327
rect 16681 7293 16715 7327
rect 16957 7293 16991 7327
rect 21281 7293 21315 7327
rect 21833 7293 21867 7327
rect 22753 7293 22787 7327
rect 27537 7293 27571 7327
rect 28273 7293 28307 7327
rect 18337 7225 18371 7259
rect 23857 7225 23891 7259
rect 15393 7157 15427 7191
rect 18153 7157 18187 7191
rect 19073 7157 19107 7191
rect 20637 7157 20671 7191
rect 23213 7157 23247 7191
rect 24823 7157 24857 7191
rect 25053 7157 25087 7191
rect 26985 7157 27019 7191
rect 30021 7157 30055 7191
rect 37657 7157 37691 7191
rect 2237 6953 2271 6987
rect 22477 6953 22511 6987
rect 27951 6953 27985 6987
rect 18613 6885 18647 6919
rect 21925 6885 21959 6919
rect 14565 6817 14599 6851
rect 16313 6817 16347 6851
rect 17141 6817 17175 6851
rect 18245 6817 18279 6851
rect 22293 6817 22327 6851
rect 25513 6817 25547 6851
rect 27721 6817 27755 6851
rect 29653 6817 29687 6851
rect 36277 6817 36311 6851
rect 37197 6817 37231 6851
rect 1685 6749 1719 6783
rect 2329 6749 2363 6783
rect 2973 6749 3007 6783
rect 16957 6749 16991 6783
rect 17233 6749 17267 6783
rect 19441 6749 19475 6783
rect 20913 6749 20947 6783
rect 21097 6749 21131 6783
rect 21373 6749 21407 6783
rect 22109 6749 22143 6783
rect 22569 6749 22603 6783
rect 23029 6749 23063 6783
rect 23397 6749 23431 6783
rect 25421 6749 25455 6783
rect 26157 6749 26191 6783
rect 26341 6749 26375 6783
rect 26801 6749 26835 6783
rect 26985 6749 27019 6783
rect 29745 6749 29779 6783
rect 14841 6681 14875 6715
rect 21005 6681 21039 6715
rect 21215 6681 21249 6715
rect 23305 6681 23339 6715
rect 25329 6681 25363 6715
rect 26249 6681 26283 6715
rect 36461 6681 36495 6715
rect 2881 6613 2915 6647
rect 16773 6613 16807 6647
rect 18705 6613 18739 6647
rect 19671 6613 19705 6647
rect 20729 6613 20763 6647
rect 23029 6613 23063 6647
rect 23213 6613 23247 6647
rect 24961 6613 24995 6647
rect 26893 6613 26927 6647
rect 15117 6409 15151 6443
rect 17065 6409 17099 6443
rect 21005 6409 21039 6443
rect 24041 6409 24075 6443
rect 25053 6409 25087 6443
rect 25513 6409 25547 6443
rect 27077 6409 27111 6443
rect 1869 6341 1903 6375
rect 16865 6341 16899 6375
rect 20453 6341 20487 6375
rect 22201 6341 22235 6375
rect 23121 6341 23155 6375
rect 28549 6341 28583 6375
rect 37657 6341 37691 6375
rect 1685 6273 1719 6307
rect 15301 6273 15335 6307
rect 17693 6273 17727 6307
rect 17877 6273 17911 6307
rect 17969 6273 18003 6307
rect 18061 6273 18095 6307
rect 18981 6273 19015 6307
rect 21005 6273 21039 6307
rect 21189 6273 21223 6307
rect 21833 6273 21867 6307
rect 22017 6273 22051 6307
rect 22845 6273 22879 6307
rect 23029 6273 23063 6307
rect 23213 6273 23247 6307
rect 23857 6273 23891 6307
rect 24133 6273 24167 6307
rect 24869 6273 24903 6307
rect 25513 6273 25547 6307
rect 25697 6273 25731 6307
rect 28825 6273 28859 6307
rect 38025 6273 38059 6307
rect 2789 6205 2823 6239
rect 18705 6205 18739 6239
rect 19993 6205 20027 6239
rect 17233 6137 17267 6171
rect 20085 6137 20119 6171
rect 17049 6069 17083 6103
rect 18245 6069 18279 6103
rect 23397 6069 23431 6103
rect 23857 6069 23891 6103
rect 36737 6069 36771 6103
rect 15485 5865 15519 5899
rect 16681 5865 16715 5899
rect 17693 5865 17727 5899
rect 19441 5865 19475 5899
rect 22109 5865 22143 5899
rect 27721 5865 27755 5899
rect 18613 5729 18647 5763
rect 20637 5729 20671 5763
rect 23305 5729 23339 5763
rect 37105 5729 37139 5763
rect 1961 5661 1995 5695
rect 2605 5661 2639 5695
rect 3249 5661 3283 5695
rect 3801 5661 3835 5695
rect 5089 5661 5123 5695
rect 15577 5661 15611 5695
rect 16037 5661 16071 5695
rect 16865 5661 16899 5695
rect 17509 5661 17543 5695
rect 17785 5661 17819 5695
rect 18521 5661 18555 5695
rect 19257 5661 19291 5695
rect 20361 5661 20395 5695
rect 23029 5661 23063 5695
rect 24409 5661 24443 5695
rect 24593 5661 24627 5695
rect 25237 5661 25271 5695
rect 25881 5661 25915 5695
rect 27813 5661 27847 5695
rect 35633 5661 35667 5695
rect 38117 5661 38151 5695
rect 1869 5593 1903 5627
rect 19349 5593 19383 5627
rect 19533 5593 19567 5627
rect 37933 5593 37967 5627
rect 2513 5525 2547 5559
rect 16129 5525 16163 5559
rect 17325 5525 17359 5559
rect 24777 5525 24811 5559
rect 25329 5525 25363 5559
rect 25973 5525 26007 5559
rect 15945 5321 15979 5355
rect 18613 5321 18647 5355
rect 20821 5321 20855 5355
rect 22937 5321 22971 5355
rect 23765 5321 23799 5355
rect 23933 5321 23967 5355
rect 24685 5321 24719 5355
rect 36645 5321 36679 5355
rect 37565 5321 37599 5355
rect 3433 5253 3467 5287
rect 17141 5253 17175 5287
rect 23029 5253 23063 5287
rect 24133 5253 24167 5287
rect 26157 5253 26191 5287
rect 3617 5185 3651 5219
rect 5365 5185 5399 5219
rect 16129 5185 16163 5219
rect 22109 5185 22143 5219
rect 36737 5185 36771 5219
rect 37473 5185 37507 5219
rect 1777 5117 1811 5151
rect 16865 5117 16899 5151
rect 19073 5117 19107 5151
rect 19349 5117 19383 5151
rect 23213 5117 23247 5151
rect 26433 5117 26467 5151
rect 4077 4981 4111 5015
rect 5273 4981 5307 5015
rect 6377 4981 6411 5015
rect 21925 4981 21959 5015
rect 22569 4981 22603 5015
rect 23949 4981 23983 5015
rect 32965 4981 32999 5015
rect 34989 4981 35023 5015
rect 36093 4981 36127 5015
rect 15564 4777 15598 4811
rect 17049 4777 17083 4811
rect 17877 4777 17911 4811
rect 21189 4777 21223 4811
rect 23581 4777 23615 4811
rect 25053 4709 25087 4743
rect 3065 4641 3099 4675
rect 3249 4641 3283 4675
rect 4997 4641 5031 4675
rect 5181 4641 5215 4675
rect 5825 4641 5859 4675
rect 9965 4641 9999 4675
rect 15301 4641 15335 4675
rect 19441 4641 19475 4675
rect 21833 4641 21867 4675
rect 26801 4641 26835 4675
rect 33149 4641 33183 4675
rect 35725 4641 35759 4675
rect 3985 4573 4019 4607
rect 7481 4573 7515 4607
rect 8309 4573 8343 4607
rect 9137 4573 9171 4607
rect 10517 4573 10551 4607
rect 17785 4573 17819 4607
rect 18521 4573 18555 4607
rect 24593 4573 24627 4607
rect 32229 4573 32263 4607
rect 35081 4573 35115 4607
rect 1409 4505 1443 4539
rect 19717 4505 19751 4539
rect 22109 4505 22143 4539
rect 26525 4505 26559 4539
rect 32413 4505 32447 4539
rect 35173 4505 35207 4539
rect 35909 4505 35943 4539
rect 37565 4505 37599 4539
rect 3893 4437 3927 4471
rect 10609 4437 10643 4471
rect 18613 4437 18647 4471
rect 24501 4437 24535 4471
rect 19901 4233 19935 4267
rect 22201 4233 22235 4267
rect 5181 4097 5215 4131
rect 7481 4097 7515 4131
rect 9965 4097 9999 4131
rect 10609 4097 10643 4131
rect 19441 4097 19475 4131
rect 20085 4097 20119 4131
rect 20729 4097 20763 4131
rect 22385 4097 22419 4131
rect 24777 4097 24811 4131
rect 25697 4097 25731 4131
rect 25789 4097 25823 4131
rect 31033 4097 31067 4131
rect 32597 4097 32631 4131
rect 36737 4097 36771 4131
rect 37289 4097 37323 4131
rect 38117 4097 38151 4131
rect 2605 4029 2639 4063
rect 4169 4029 4203 4063
rect 4353 4029 4387 4063
rect 7665 4029 7699 4063
rect 8861 4029 8895 4063
rect 23029 4029 23063 4063
rect 24501 4029 24535 4063
rect 32781 4029 32815 4063
rect 33517 4029 33551 4063
rect 35817 4029 35851 4063
rect 36553 4029 36587 4063
rect 2053 3961 2087 3995
rect 5089 3961 5123 3995
rect 19349 3961 19383 3995
rect 5825 3893 5859 3927
rect 6377 3893 6411 3927
rect 9873 3893 9907 3927
rect 10517 3893 10551 3927
rect 11529 3893 11563 3927
rect 13277 3893 13311 3927
rect 20821 3893 20855 3927
rect 31125 3893 31159 3927
rect 8309 3689 8343 3723
rect 23121 3689 23155 3723
rect 33425 3689 33459 3723
rect 37841 3689 37875 3723
rect 4721 3553 4755 3587
rect 5917 3553 5951 3587
rect 8953 3553 8987 3587
rect 10609 3553 10643 3587
rect 10793 3553 10827 3587
rect 11253 3553 11287 3587
rect 11437 3553 11471 3587
rect 11713 3553 11747 3587
rect 15117 3553 15151 3587
rect 21189 3553 21223 3587
rect 22385 3553 22419 3587
rect 31217 3553 31251 3587
rect 31585 3553 31619 3587
rect 35449 3553 35483 3587
rect 36829 3553 36863 3587
rect 1685 3485 1719 3519
rect 2329 3485 2363 3519
rect 2789 3485 2823 3519
rect 6377 3485 6411 3519
rect 7573 3485 7607 3519
rect 8401 3485 8435 3519
rect 14657 3485 14691 3519
rect 16313 3485 16347 3519
rect 17601 3485 17635 3519
rect 18429 3485 18463 3519
rect 19717 3485 19751 3519
rect 22569 3485 22603 3519
rect 23213 3485 23247 3519
rect 24685 3485 24719 3519
rect 30573 3485 30607 3519
rect 31033 3485 31067 3519
rect 33517 3485 33551 3519
rect 33977 3485 34011 3519
rect 34805 3485 34839 3519
rect 37749 3485 37783 3519
rect 5733 3417 5767 3451
rect 34897 3417 34931 3451
rect 35633 3417 35667 3451
rect 2237 3349 2271 3383
rect 2881 3349 2915 3383
rect 7665 3349 7699 3383
rect 14565 3349 14599 3383
rect 16405 3349 16439 3383
rect 17693 3349 17727 3383
rect 19625 3349 19659 3383
rect 24777 3349 24811 3383
rect 34069 3349 34103 3383
rect 4353 3145 4387 3179
rect 30849 3145 30883 3179
rect 1961 3077 1995 3111
rect 5733 3077 5767 3111
rect 6561 3077 6595 3111
rect 9229 3077 9263 3111
rect 14473 3077 14507 3111
rect 16865 3077 16899 3111
rect 19165 3077 19199 3111
rect 24777 3077 24811 3111
rect 31493 3077 31527 3111
rect 32321 3077 32355 3111
rect 35081 3077 35115 3111
rect 1777 3009 1811 3043
rect 4445 3009 4479 3043
rect 5089 3009 5123 3043
rect 5641 3009 5675 3043
rect 6377 3009 6411 3043
rect 9045 3009 9079 3043
rect 13829 3009 13863 3043
rect 14289 3009 14323 3043
rect 18981 3009 19015 3043
rect 30757 3009 30791 3043
rect 31401 3009 31435 3043
rect 34897 3009 34931 3043
rect 37381 3009 37415 3043
rect 2789 2941 2823 2975
rect 6837 2941 6871 2975
rect 9689 2941 9723 2975
rect 13369 2941 13403 2975
rect 13645 2941 13679 2975
rect 14841 2941 14875 2975
rect 16681 2941 16715 2975
rect 17141 2941 17175 2975
rect 19441 2941 19475 2975
rect 21833 2941 21867 2975
rect 22017 2941 22051 2975
rect 22569 2941 22603 2975
rect 24593 2941 24627 2975
rect 25145 2941 25179 2975
rect 32137 2941 32171 2975
rect 32597 2941 32631 2975
rect 35449 2941 35483 2975
rect 4997 2805 5031 2839
rect 37473 2805 37507 2839
rect 13277 2601 13311 2635
rect 16681 2601 16715 2635
rect 21925 2601 21959 2635
rect 22477 2601 22511 2635
rect 23121 2601 23155 2635
rect 24685 2601 24719 2635
rect 31585 2601 31619 2635
rect 37933 2601 37967 2635
rect 30941 2533 30975 2567
rect 37381 2533 37415 2567
rect 3065 2465 3099 2499
rect 3249 2465 3283 2499
rect 5457 2465 5491 2499
rect 5641 2465 5675 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 9413 2465 9447 2499
rect 19533 2465 19567 2499
rect 19993 2465 20027 2499
rect 33701 2465 33735 2499
rect 33977 2465 34011 2499
rect 36553 2465 36587 2499
rect 36737 2465 36771 2499
rect 8953 2397 8987 2431
rect 13369 2397 13403 2431
rect 18705 2397 18739 2431
rect 19349 2397 19383 2431
rect 21833 2397 21867 2431
rect 34161 2397 34195 2431
rect 37289 2397 37323 2431
rect 1409 2329 1443 2363
rect 3801 2329 3835 2363
rect 9137 2329 9171 2363
rect 34897 2329 34931 2363
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 10597 37383 10655 37389
rect 10597 37349 10609 37383
rect 10643 37380 10655 37383
rect 11514 37380 11520 37392
rect 10643 37352 11520 37380
rect 10643 37349 10655 37352
rect 10597 37343 10655 37349
rect 11514 37340 11520 37352
rect 11572 37340 11578 37392
rect 34149 37383 34207 37389
rect 34149 37349 34161 37383
rect 34195 37380 34207 37383
rect 34882 37380 34888 37392
rect 34195 37352 34888 37380
rect 34195 37349 34207 37352
rect 34149 37343 34207 37349
rect 34882 37340 34888 37352
rect 34940 37340 34946 37392
rect 9309 37315 9367 37321
rect 9309 37281 9321 37315
rect 9355 37312 9367 37315
rect 9355 37284 11560 37312
rect 9355 37281 9367 37284
rect 9309 37275 9367 37281
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 2130 37204 2136 37256
rect 2188 37244 2194 37256
rect 2317 37247 2375 37253
rect 2317 37244 2329 37247
rect 2188 37216 2329 37244
rect 2188 37204 2194 37216
rect 2317 37213 2329 37216
rect 2363 37213 2375 37247
rect 2317 37207 2375 37213
rect 2961 37247 3019 37253
rect 2961 37213 2973 37247
rect 3007 37244 3019 37247
rect 3007 37216 4292 37244
rect 3007 37213 3019 37216
rect 2961 37207 3019 37213
rect 1946 37136 1952 37188
rect 2004 37176 2010 37188
rect 3789 37179 3847 37185
rect 3789 37176 3801 37179
rect 2004 37148 3801 37176
rect 2004 37136 2010 37148
rect 3789 37145 3801 37148
rect 3835 37145 3847 37179
rect 3789 37139 3847 37145
rect 1581 37111 1639 37117
rect 1581 37077 1593 37111
rect 1627 37108 1639 37111
rect 2038 37108 2044 37120
rect 1627 37080 2044 37108
rect 1627 37077 1639 37080
rect 1581 37071 1639 37077
rect 2038 37068 2044 37080
rect 2096 37068 2102 37120
rect 2222 37108 2228 37120
rect 2183 37080 2228 37108
rect 2222 37068 2228 37080
rect 2280 37068 2286 37120
rect 2869 37111 2927 37117
rect 2869 37077 2881 37111
rect 2915 37108 2927 37111
rect 3050 37108 3056 37120
rect 2915 37080 3056 37108
rect 2915 37077 2927 37080
rect 2869 37071 2927 37077
rect 3050 37068 3056 37080
rect 3108 37068 3114 37120
rect 4264 37108 4292 37216
rect 5626 37204 5632 37256
rect 5684 37244 5690 37256
rect 6638 37244 6644 37256
rect 5684 37216 5729 37244
rect 6599 37216 6644 37244
rect 5684 37204 5690 37216
rect 6638 37204 6644 37216
rect 6696 37204 6702 37256
rect 7285 37247 7343 37253
rect 7285 37213 7297 37247
rect 7331 37213 7343 37247
rect 7742 37244 7748 37256
rect 7703 37216 7748 37244
rect 7285 37207 7343 37213
rect 5445 37179 5503 37185
rect 5445 37145 5457 37179
rect 5491 37176 5503 37179
rect 7193 37179 7251 37185
rect 7193 37176 7205 37179
rect 5491 37148 7205 37176
rect 5491 37145 5503 37148
rect 5445 37139 5503 37145
rect 7193 37145 7205 37148
rect 7239 37145 7251 37179
rect 7193 37139 7251 37145
rect 7300 37120 7328 37207
rect 7742 37204 7748 37216
rect 7800 37204 7806 37256
rect 9766 37244 9772 37256
rect 9727 37216 9772 37244
rect 9766 37204 9772 37216
rect 9824 37204 9830 37256
rect 11532 37253 11560 37284
rect 11698 37272 11704 37324
rect 11756 37312 11762 37324
rect 11977 37315 12035 37321
rect 11977 37312 11989 37315
rect 11756 37284 11989 37312
rect 11756 37272 11762 37284
rect 11977 37281 11989 37284
rect 12023 37281 12035 37315
rect 11977 37275 12035 37281
rect 14921 37315 14979 37321
rect 14921 37281 14933 37315
rect 14967 37312 14979 37315
rect 16114 37312 16120 37324
rect 14967 37284 16120 37312
rect 14967 37281 14979 37284
rect 14921 37275 14979 37281
rect 16114 37272 16120 37284
rect 16172 37272 16178 37324
rect 17221 37315 17279 37321
rect 17221 37281 17233 37315
rect 17267 37312 17279 37315
rect 20622 37312 20628 37324
rect 17267 37284 19472 37312
rect 20583 37284 20628 37312
rect 17267 37281 17279 37284
rect 17221 37275 17279 37281
rect 11517 37247 11575 37253
rect 11517 37213 11529 37247
rect 11563 37213 11575 37247
rect 11517 37207 11575 37213
rect 14093 37247 14151 37253
rect 14093 37213 14105 37247
rect 14139 37213 14151 37247
rect 17678 37244 17684 37256
rect 17639 37216 17684 37244
rect 14093 37207 14151 37213
rect 10870 37136 10876 37188
rect 10928 37176 10934 37188
rect 11701 37179 11759 37185
rect 11701 37176 11713 37179
rect 10928 37148 11713 37176
rect 10928 37136 10934 37148
rect 11701 37145 11713 37148
rect 11747 37145 11759 37179
rect 11701 37139 11759 37145
rect 12158 37136 12164 37188
rect 12216 37176 12222 37188
rect 14108 37176 14136 37207
rect 17678 37204 17684 37216
rect 17736 37204 17742 37256
rect 18690 37244 18696 37256
rect 18651 37216 18696 37244
rect 18690 37204 18696 37216
rect 18748 37204 18754 37256
rect 19444 37253 19472 37284
rect 20622 37272 20628 37284
rect 20680 37272 20686 37324
rect 27246 37312 27252 37324
rect 27207 37284 27252 37312
rect 27246 37272 27252 37284
rect 27304 37272 27310 37324
rect 32125 37315 32183 37321
rect 32125 37312 32137 37315
rect 29748 37284 32137 37312
rect 19429 37247 19487 37253
rect 19429 37213 19441 37247
rect 19475 37213 19487 37247
rect 21818 37244 21824 37256
rect 21779 37216 21824 37244
rect 19429 37207 19487 37213
rect 21818 37204 21824 37216
rect 21876 37204 21882 37256
rect 23017 37247 23075 37253
rect 23017 37213 23029 37247
rect 23063 37244 23075 37247
rect 23106 37244 23112 37256
rect 23063 37216 23112 37244
rect 23063 37213 23075 37216
rect 23017 37207 23075 37213
rect 23106 37204 23112 37216
rect 23164 37204 23170 37256
rect 23658 37244 23664 37256
rect 23619 37216 23664 37244
rect 23658 37204 23664 37216
rect 23716 37204 23722 37256
rect 24118 37204 24124 37256
rect 24176 37244 24182 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 24176 37216 24409 37244
rect 24176 37204 24182 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 25406 37244 25412 37256
rect 25367 37216 25412 37244
rect 24397 37207 24455 37213
rect 25406 37204 25412 37216
rect 25464 37204 25470 37256
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25832 37216 25881 37244
rect 25832 37204 25838 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 26142 37204 26148 37256
rect 26200 37244 26206 37256
rect 29748 37253 29776 37284
rect 32125 37281 32137 37284
rect 32171 37281 32183 37315
rect 32125 37275 32183 37281
rect 33505 37315 33563 37321
rect 33505 37281 33517 37315
rect 33551 37312 33563 37315
rect 36722 37312 36728 37324
rect 33551 37284 34928 37312
rect 36683 37284 36728 37312
rect 33551 37281 33563 37284
rect 33505 37275 33563 37281
rect 34900 37253 34928 37284
rect 36722 37272 36728 37284
rect 36780 37272 36786 37324
rect 26973 37247 27031 37253
rect 26973 37244 26985 37247
rect 26200 37216 26985 37244
rect 26200 37204 26206 37216
rect 26973 37213 26985 37216
rect 27019 37213 27031 37247
rect 26973 37207 27031 37213
rect 29733 37247 29791 37253
rect 29733 37213 29745 37247
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 34885 37247 34943 37253
rect 34885 37213 34897 37247
rect 34931 37213 34943 37247
rect 37274 37244 37280 37256
rect 37235 37216 37280 37244
rect 34885 37207 34943 37213
rect 37274 37204 37280 37216
rect 37332 37204 37338 37256
rect 37918 37244 37924 37256
rect 37879 37216 37924 37244
rect 37918 37204 37924 37216
rect 37976 37204 37982 37256
rect 12216 37148 14136 37176
rect 19613 37179 19671 37185
rect 12216 37136 12222 37148
rect 19613 37145 19625 37179
rect 19659 37176 19671 37179
rect 19659 37148 19748 37176
rect 19659 37145 19671 37148
rect 19613 37139 19671 37145
rect 19720 37147 19748 37148
rect 5810 37108 5816 37120
rect 4264 37080 5816 37108
rect 5810 37068 5816 37080
rect 5868 37068 5874 37120
rect 6454 37108 6460 37120
rect 6415 37080 6460 37108
rect 6454 37068 6460 37080
rect 6512 37068 6518 37120
rect 7282 37108 7288 37120
rect 7195 37080 7288 37108
rect 7282 37068 7288 37080
rect 7340 37108 7346 37120
rect 12710 37108 12716 37120
rect 7340 37080 12716 37108
rect 7340 37068 7346 37080
rect 12710 37068 12716 37080
rect 12768 37068 12774 37120
rect 14182 37108 14188 37120
rect 14143 37080 14188 37108
rect 14182 37068 14188 37080
rect 14240 37068 14246 37120
rect 19720 37119 19840 37147
rect 20070 37136 20076 37188
rect 20128 37176 20134 37188
rect 22370 37176 22376 37188
rect 20128 37148 22376 37176
rect 20128 37136 20134 37148
rect 22370 37136 22376 37148
rect 22428 37136 22434 37188
rect 29546 37176 29552 37188
rect 28474 37148 29552 37176
rect 29546 37136 29552 37148
rect 29604 37136 29610 37188
rect 29638 37136 29644 37188
rect 29696 37176 29702 37188
rect 29917 37179 29975 37185
rect 29917 37176 29929 37179
rect 29696 37148 29929 37176
rect 29696 37136 29702 37148
rect 29917 37145 29929 37148
rect 29963 37145 29975 37179
rect 29917 37139 29975 37145
rect 30926 37136 30932 37188
rect 30984 37176 30990 37188
rect 31573 37179 31631 37185
rect 31573 37176 31585 37179
rect 30984 37148 31585 37176
rect 30984 37136 30990 37148
rect 31573 37145 31585 37148
rect 31619 37145 31631 37179
rect 31573 37139 31631 37145
rect 34790 37136 34796 37188
rect 34848 37176 34854 37188
rect 35069 37179 35127 37185
rect 35069 37176 35081 37179
rect 34848 37148 35081 37176
rect 34848 37136 34854 37148
rect 35069 37145 35081 37148
rect 35115 37145 35127 37179
rect 35069 37139 35127 37145
rect 36538 37136 36544 37188
rect 36596 37176 36602 37188
rect 38013 37179 38071 37185
rect 38013 37176 38025 37179
rect 36596 37148 38025 37176
rect 36596 37136 36602 37148
rect 38013 37145 38025 37148
rect 38059 37145 38071 37179
rect 38013 37139 38071 37145
rect 19812 37108 19840 37119
rect 21726 37108 21732 37120
rect 19812 37080 21732 37108
rect 21726 37068 21732 37080
rect 21784 37068 21790 37120
rect 21910 37108 21916 37120
rect 21871 37080 21916 37108
rect 21910 37068 21916 37080
rect 21968 37068 21974 37120
rect 22830 37068 22836 37120
rect 22888 37108 22894 37120
rect 22925 37111 22983 37117
rect 22925 37108 22937 37111
rect 22888 37080 22937 37108
rect 22888 37068 22894 37080
rect 22925 37077 22937 37080
rect 22971 37077 22983 37111
rect 25958 37108 25964 37120
rect 25919 37080 25964 37108
rect 22925 37071 22983 37077
rect 25958 37068 25964 37080
rect 26016 37068 26022 37120
rect 28718 37108 28724 37120
rect 28679 37080 28724 37108
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 35894 37068 35900 37120
rect 35952 37108 35958 37120
rect 37369 37111 37427 37117
rect 37369 37108 37381 37111
rect 35952 37080 37381 37108
rect 35952 37068 35958 37080
rect 37369 37077 37381 37080
rect 37415 37077 37427 37111
rect 37369 37071 37427 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 2038 36864 2044 36916
rect 2096 36904 2102 36916
rect 5718 36904 5724 36916
rect 2096 36876 5724 36904
rect 2096 36864 2102 36876
rect 5718 36864 5724 36876
rect 5776 36904 5782 36916
rect 6638 36904 6644 36916
rect 5776 36876 6644 36904
rect 5776 36864 5782 36876
rect 6638 36864 6644 36876
rect 6696 36864 6702 36916
rect 10870 36904 10876 36916
rect 10831 36876 10876 36904
rect 10870 36864 10876 36876
rect 10928 36864 10934 36916
rect 12618 36904 12624 36916
rect 10980 36876 12624 36904
rect 1578 36836 1584 36848
rect 1539 36808 1584 36836
rect 1578 36796 1584 36808
rect 1636 36796 1642 36848
rect 2222 36796 2228 36848
rect 2280 36836 2286 36848
rect 3237 36839 3295 36845
rect 3237 36836 3249 36839
rect 2280 36808 3249 36836
rect 2280 36796 2286 36808
rect 3237 36805 3249 36808
rect 3283 36805 3295 36839
rect 3878 36836 3884 36848
rect 3839 36808 3884 36836
rect 3237 36799 3295 36805
rect 3878 36796 3884 36808
rect 3936 36796 3942 36848
rect 7742 36836 7748 36848
rect 5736 36808 7748 36836
rect 5736 36777 5764 36808
rect 7742 36796 7748 36808
rect 7800 36796 7806 36848
rect 10502 36796 10508 36848
rect 10560 36836 10566 36848
rect 10980 36836 11008 36876
rect 12618 36864 12624 36876
rect 12676 36864 12682 36916
rect 12710 36864 12716 36916
rect 12768 36904 12774 36916
rect 23106 36904 23112 36916
rect 12768 36876 23112 36904
rect 12768 36864 12774 36876
rect 23106 36864 23112 36876
rect 23164 36864 23170 36916
rect 25774 36864 25780 36916
rect 25832 36904 25838 36916
rect 25832 36876 37596 36904
rect 25832 36864 25838 36876
rect 12066 36836 12072 36848
rect 10560 36808 11008 36836
rect 11072 36808 12072 36836
rect 10560 36796 10566 36808
rect 5721 36771 5779 36777
rect 5721 36737 5733 36771
rect 5767 36737 5779 36771
rect 6454 36768 6460 36780
rect 6415 36740 6460 36768
rect 5721 36731 5779 36737
rect 6454 36728 6460 36740
rect 6512 36728 6518 36780
rect 7190 36768 7196 36780
rect 7151 36740 7196 36768
rect 7190 36728 7196 36740
rect 7248 36728 7254 36780
rect 10410 36728 10416 36780
rect 10468 36768 10474 36780
rect 10781 36771 10839 36777
rect 10781 36768 10793 36771
rect 10468 36740 10793 36768
rect 10468 36728 10474 36740
rect 10781 36737 10793 36740
rect 10827 36768 10839 36771
rect 11072 36768 11100 36808
rect 12066 36796 12072 36808
rect 12124 36796 12130 36848
rect 12250 36796 12256 36848
rect 12308 36836 12314 36848
rect 14277 36839 14335 36845
rect 14277 36836 14289 36839
rect 12308 36808 14289 36836
rect 12308 36796 12314 36808
rect 14277 36805 14289 36808
rect 14323 36805 14335 36839
rect 14277 36799 14335 36805
rect 14752 36808 20852 36836
rect 11514 36768 11520 36780
rect 10827 36740 11100 36768
rect 11475 36740 11520 36768
rect 10827 36737 10839 36740
rect 10781 36731 10839 36737
rect 11514 36728 11520 36740
rect 11572 36728 11578 36780
rect 3418 36700 3424 36712
rect 3379 36672 3424 36700
rect 3418 36660 3424 36672
rect 3476 36660 3482 36712
rect 5534 36700 5540 36712
rect 5495 36672 5540 36700
rect 5534 36660 5540 36672
rect 5592 36660 5598 36712
rect 8386 36700 8392 36712
rect 8347 36672 8392 36700
rect 8386 36660 8392 36672
rect 8444 36660 8450 36712
rect 8573 36703 8631 36709
rect 8573 36669 8585 36703
rect 8619 36700 8631 36703
rect 9030 36700 9036 36712
rect 8619 36672 9036 36700
rect 8619 36669 8631 36672
rect 8573 36663 8631 36669
rect 9030 36660 9036 36672
rect 9088 36660 9094 36712
rect 9769 36703 9827 36709
rect 9769 36700 9781 36703
rect 9692 36672 9781 36700
rect 9692 36644 9720 36672
rect 9769 36669 9781 36672
rect 9815 36669 9827 36703
rect 11698 36700 11704 36712
rect 11659 36672 11704 36700
rect 9769 36663 9827 36669
rect 11698 36660 11704 36672
rect 11756 36660 11762 36712
rect 11977 36703 12035 36709
rect 11977 36669 11989 36703
rect 12023 36669 12035 36703
rect 11977 36663 12035 36669
rect 9674 36592 9680 36644
rect 9732 36592 9738 36644
rect 10962 36592 10968 36644
rect 11020 36632 11026 36644
rect 11992 36632 12020 36663
rect 12066 36660 12072 36712
rect 12124 36700 12130 36712
rect 14752 36700 14780 36808
rect 16114 36728 16120 36780
rect 16172 36768 16178 36780
rect 17126 36768 17132 36780
rect 16172 36740 16217 36768
rect 17087 36740 17132 36768
rect 16172 36728 16178 36740
rect 17126 36728 17132 36740
rect 17184 36728 17190 36780
rect 17678 36768 17684 36780
rect 17639 36740 17684 36768
rect 17678 36728 17684 36740
rect 17736 36728 17742 36780
rect 12124 36672 14780 36700
rect 15933 36703 15991 36709
rect 12124 36660 12130 36672
rect 15933 36669 15945 36703
rect 15979 36700 15991 36703
rect 17034 36700 17040 36712
rect 15979 36672 17040 36700
rect 15979 36669 15991 36672
rect 15933 36663 15991 36669
rect 17034 36660 17040 36672
rect 17092 36660 17098 36712
rect 17862 36700 17868 36712
rect 17823 36672 17868 36700
rect 17862 36660 17868 36672
rect 17920 36660 17926 36712
rect 18046 36660 18052 36712
rect 18104 36700 18110 36712
rect 18141 36703 18199 36709
rect 18141 36700 18153 36703
rect 18104 36672 18153 36700
rect 18104 36660 18110 36672
rect 18141 36669 18153 36672
rect 18187 36669 18199 36703
rect 18141 36663 18199 36669
rect 20717 36703 20775 36709
rect 20717 36669 20729 36703
rect 20763 36669 20775 36703
rect 20824 36700 20852 36808
rect 21266 36796 21272 36848
rect 21324 36836 21330 36848
rect 21821 36839 21879 36845
rect 21821 36836 21833 36839
rect 21324 36808 21833 36836
rect 21324 36796 21330 36808
rect 21821 36805 21833 36808
rect 21867 36805 21879 36839
rect 28537 36839 28595 36845
rect 21821 36799 21879 36805
rect 22066 36808 27844 36836
rect 21174 36768 21180 36780
rect 21135 36740 21180 36768
rect 21174 36728 21180 36740
rect 21232 36728 21238 36780
rect 22066 36768 22094 36808
rect 21284 36740 22094 36768
rect 21284 36700 21312 36740
rect 23658 36728 23664 36780
rect 23716 36768 23722 36780
rect 24118 36768 24124 36780
rect 23716 36740 23761 36768
rect 24079 36740 24124 36768
rect 23716 36728 23722 36740
rect 24118 36728 24124 36740
rect 24176 36728 24182 36780
rect 27816 36777 27844 36808
rect 28537 36805 28549 36839
rect 28583 36836 28595 36839
rect 29273 36839 29331 36845
rect 29273 36836 29285 36839
rect 28583 36808 29285 36836
rect 28583 36805 28595 36808
rect 28537 36799 28595 36805
rect 29273 36805 29285 36808
rect 29319 36805 29331 36839
rect 29273 36799 29331 36805
rect 35069 36839 35127 36845
rect 35069 36805 35081 36839
rect 35115 36836 35127 36839
rect 37461 36839 37519 36845
rect 37461 36836 37473 36839
rect 35115 36808 37473 36836
rect 35115 36805 35127 36808
rect 35069 36799 35127 36805
rect 37461 36805 37473 36808
rect 37507 36805 37519 36839
rect 37461 36799 37519 36805
rect 27801 36771 27859 36777
rect 27801 36737 27813 36771
rect 27847 36768 27859 36771
rect 28258 36768 28264 36780
rect 27847 36740 28264 36768
rect 27847 36737 27859 36740
rect 27801 36731 27859 36737
rect 28258 36728 28264 36740
rect 28316 36728 28322 36780
rect 28445 36771 28503 36777
rect 28445 36737 28457 36771
rect 28491 36737 28503 36771
rect 34882 36768 34888 36780
rect 34843 36740 34888 36768
rect 28445 36731 28503 36737
rect 20824 36672 21312 36700
rect 20717 36663 20775 36669
rect 20732 36632 20760 36663
rect 21910 36660 21916 36712
rect 21968 36700 21974 36712
rect 23477 36703 23535 36709
rect 23477 36700 23489 36703
rect 21968 36672 23489 36700
rect 21968 36660 21974 36672
rect 23477 36669 23489 36672
rect 23523 36669 23535 36703
rect 23477 36663 23535 36669
rect 24305 36703 24363 36709
rect 24305 36669 24317 36703
rect 24351 36700 24363 36703
rect 24486 36700 24492 36712
rect 24351 36672 24492 36700
rect 24351 36669 24363 36672
rect 24305 36663 24363 36669
rect 24486 36660 24492 36672
rect 24544 36660 24550 36712
rect 24578 36660 24584 36712
rect 24636 36700 24642 36712
rect 28460 36700 28488 36731
rect 34882 36728 34888 36740
rect 34940 36728 34946 36780
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36768 36783 36771
rect 37182 36768 37188 36780
rect 36771 36740 37188 36768
rect 36771 36737 36783 36740
rect 36725 36731 36783 36737
rect 37182 36728 37188 36740
rect 37240 36728 37246 36780
rect 37369 36771 37427 36777
rect 37369 36737 37381 36771
rect 37415 36768 37427 36771
rect 37568 36768 37596 36876
rect 38562 36768 38568 36780
rect 37415 36740 38568 36768
rect 37415 36737 37427 36740
rect 37369 36731 37427 36737
rect 38562 36728 38568 36740
rect 38620 36728 38626 36780
rect 28994 36700 29000 36712
rect 24636 36672 24681 36700
rect 27264 36672 29000 36700
rect 24636 36660 24642 36672
rect 26786 36632 26792 36644
rect 11020 36604 12020 36632
rect 16868 36604 26792 36632
rect 11020 36592 11026 36604
rect 10686 36524 10692 36576
rect 10744 36564 10750 36576
rect 16868 36564 16896 36604
rect 26786 36592 26792 36604
rect 26844 36592 26850 36644
rect 10744 36536 16896 36564
rect 10744 36524 10750 36536
rect 16942 36524 16948 36576
rect 17000 36564 17006 36576
rect 17037 36567 17095 36573
rect 17037 36564 17049 36567
rect 17000 36536 17049 36564
rect 17000 36524 17006 36536
rect 17037 36533 17049 36536
rect 17083 36533 17095 36567
rect 17037 36527 17095 36533
rect 17126 36524 17132 36576
rect 17184 36564 17190 36576
rect 19426 36564 19432 36576
rect 17184 36536 19432 36564
rect 17184 36524 17190 36536
rect 19426 36524 19432 36536
rect 19484 36524 19490 36576
rect 21634 36524 21640 36576
rect 21692 36564 21698 36576
rect 27264 36564 27292 36672
rect 28994 36660 29000 36672
rect 29052 36660 29058 36712
rect 29089 36703 29147 36709
rect 29089 36669 29101 36703
rect 29135 36700 29147 36703
rect 30190 36700 30196 36712
rect 29135 36672 30196 36700
rect 29135 36669 29147 36672
rect 29089 36663 29147 36669
rect 30190 36660 30196 36672
rect 30248 36660 30254 36712
rect 30469 36703 30527 36709
rect 30469 36669 30481 36703
rect 30515 36669 30527 36703
rect 32398 36700 32404 36712
rect 32359 36672 32404 36700
rect 30469 36663 30527 36669
rect 29730 36592 29736 36644
rect 29788 36632 29794 36644
rect 30484 36632 30512 36663
rect 32398 36660 32404 36672
rect 32456 36660 32462 36712
rect 32582 36700 32588 36712
rect 32543 36672 32588 36700
rect 32582 36660 32588 36672
rect 32640 36660 32646 36712
rect 32858 36700 32864 36712
rect 32819 36672 32864 36700
rect 32858 36660 32864 36672
rect 32916 36660 32922 36712
rect 29788 36604 30512 36632
rect 29788 36592 29794 36604
rect 21692 36536 27292 36564
rect 27341 36567 27399 36573
rect 21692 36524 21698 36536
rect 27341 36533 27353 36567
rect 27387 36564 27399 36567
rect 27798 36564 27804 36576
rect 27387 36536 27804 36564
rect 27387 36533 27399 36536
rect 27341 36527 27399 36533
rect 27798 36524 27804 36536
rect 27856 36524 27862 36576
rect 27893 36567 27951 36573
rect 27893 36533 27905 36567
rect 27939 36564 27951 36567
rect 27982 36564 27988 36576
rect 27939 36536 27988 36564
rect 27939 36533 27951 36536
rect 27893 36527 27951 36533
rect 27982 36524 27988 36536
rect 28040 36524 28046 36576
rect 31573 36567 31631 36573
rect 31573 36533 31585 36567
rect 31619 36564 31631 36567
rect 31662 36564 31668 36576
rect 31619 36536 31668 36564
rect 31619 36533 31631 36536
rect 31573 36527 31631 36533
rect 31662 36524 31668 36536
rect 31720 36524 31726 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 9030 36360 9036 36372
rect 8991 36332 9036 36360
rect 9030 36320 9036 36332
rect 9088 36320 9094 36372
rect 9858 36320 9864 36372
rect 9916 36360 9922 36372
rect 10410 36360 10416 36372
rect 9916 36332 10416 36360
rect 9916 36320 9922 36332
rect 10410 36320 10416 36332
rect 10468 36320 10474 36372
rect 12618 36320 12624 36372
rect 12676 36360 12682 36372
rect 17034 36360 17040 36372
rect 12676 36332 15792 36360
rect 16995 36332 17040 36360
rect 12676 36320 12682 36332
rect 2130 36252 2136 36304
rect 2188 36292 2194 36304
rect 15764 36292 15792 36332
rect 17034 36320 17040 36332
rect 17092 36320 17098 36372
rect 17862 36360 17868 36372
rect 17823 36332 17868 36360
rect 17862 36320 17868 36332
rect 17920 36320 17926 36372
rect 20070 36360 20076 36372
rect 17972 36332 20076 36360
rect 17972 36292 18000 36332
rect 20070 36320 20076 36332
rect 20128 36320 20134 36372
rect 24486 36360 24492 36372
rect 24447 36332 24492 36360
rect 24486 36320 24492 36332
rect 24544 36320 24550 36372
rect 29638 36360 29644 36372
rect 29599 36332 29644 36360
rect 29638 36320 29644 36332
rect 29696 36320 29702 36372
rect 30190 36360 30196 36372
rect 30151 36332 30196 36360
rect 30190 36320 30196 36332
rect 30248 36320 30254 36372
rect 34790 36360 34796 36372
rect 34751 36332 34796 36360
rect 34790 36320 34796 36332
rect 34848 36320 34854 36372
rect 2188 36264 11100 36292
rect 15764 36264 18000 36292
rect 2188 36252 2194 36264
rect 1302 36184 1308 36236
rect 1360 36224 1366 36236
rect 1397 36227 1455 36233
rect 1397 36224 1409 36227
rect 1360 36196 1409 36224
rect 1360 36184 1366 36196
rect 1397 36193 1409 36196
rect 1443 36193 1455 36227
rect 3050 36224 3056 36236
rect 3011 36196 3056 36224
rect 1397 36187 1455 36193
rect 3050 36184 3056 36196
rect 3108 36184 3114 36236
rect 4614 36224 4620 36236
rect 4575 36196 4620 36224
rect 4614 36184 4620 36196
rect 4672 36184 4678 36236
rect 5813 36227 5871 36233
rect 5813 36193 5825 36227
rect 5859 36224 5871 36227
rect 7745 36227 7803 36233
rect 7745 36224 7757 36227
rect 5859 36196 7757 36224
rect 5859 36193 5871 36196
rect 5813 36187 5871 36193
rect 7745 36193 7757 36196
rect 7791 36193 7803 36227
rect 9766 36224 9772 36236
rect 9727 36196 9772 36224
rect 7745 36187 7803 36193
rect 9766 36184 9772 36196
rect 9824 36184 9830 36236
rect 10318 36224 10324 36236
rect 10279 36196 10324 36224
rect 10318 36184 10324 36196
rect 10376 36184 10382 36236
rect 11072 36224 11100 36264
rect 18506 36252 18512 36304
rect 18564 36292 18570 36304
rect 22002 36292 22008 36304
rect 18564 36264 22008 36292
rect 18564 36252 18570 36264
rect 22002 36252 22008 36264
rect 22060 36252 22066 36304
rect 16298 36224 16304 36236
rect 11072 36196 16304 36224
rect 16298 36184 16304 36196
rect 16356 36184 16362 36236
rect 18690 36184 18696 36236
rect 18748 36224 18754 36236
rect 19245 36227 19303 36233
rect 19245 36224 19257 36227
rect 18748 36196 19257 36224
rect 18748 36184 18754 36196
rect 19245 36193 19257 36196
rect 19291 36193 19303 36227
rect 19978 36224 19984 36236
rect 19939 36196 19984 36224
rect 19245 36187 19303 36193
rect 19978 36184 19984 36196
rect 20036 36184 20042 36236
rect 25406 36184 25412 36236
rect 25464 36224 25470 36236
rect 25777 36227 25835 36233
rect 25777 36224 25789 36227
rect 25464 36196 25789 36224
rect 25464 36184 25470 36196
rect 25777 36193 25789 36196
rect 25823 36193 25835 36227
rect 25958 36224 25964 36236
rect 25919 36196 25964 36224
rect 25777 36187 25835 36193
rect 25958 36184 25964 36196
rect 26016 36184 26022 36236
rect 26418 36224 26424 36236
rect 26379 36196 26424 36224
rect 26418 36184 26424 36196
rect 26476 36184 26482 36236
rect 31662 36224 31668 36236
rect 31623 36196 31668 36224
rect 31662 36184 31668 36196
rect 31720 36184 31726 36236
rect 32214 36224 32220 36236
rect 32175 36196 32220 36224
rect 32214 36184 32220 36196
rect 32272 36184 32278 36236
rect 38102 36224 38108 36236
rect 38063 36196 38108 36224
rect 38102 36184 38108 36196
rect 38160 36184 38166 36236
rect 3237 36159 3295 36165
rect 3237 36125 3249 36159
rect 3283 36125 3295 36159
rect 6454 36156 6460 36168
rect 6415 36128 6460 36156
rect 3237 36119 3295 36125
rect 2958 36048 2964 36100
rect 3016 36088 3022 36100
rect 3252 36088 3280 36119
rect 6454 36116 6460 36128
rect 6512 36116 6518 36168
rect 8846 36116 8852 36168
rect 8904 36156 8910 36168
rect 9125 36159 9183 36165
rect 9125 36156 9137 36159
rect 8904 36128 9137 36156
rect 8904 36116 8910 36128
rect 9125 36125 9137 36128
rect 9171 36125 9183 36159
rect 12158 36156 12164 36168
rect 12119 36128 12164 36156
rect 9125 36119 9183 36125
rect 12158 36116 12164 36128
rect 12216 36116 12222 36168
rect 12989 36159 13047 36165
rect 12989 36125 13001 36159
rect 13035 36156 13047 36159
rect 13538 36156 13544 36168
rect 13035 36128 13544 36156
rect 13035 36125 13047 36128
rect 12989 36119 13047 36125
rect 13538 36116 13544 36128
rect 13596 36116 13602 36168
rect 15841 36159 15899 36165
rect 15841 36125 15853 36159
rect 15887 36156 15899 36159
rect 16390 36156 16396 36168
rect 15887 36128 16396 36156
rect 15887 36125 15899 36128
rect 15841 36119 15899 36125
rect 16390 36116 16396 36128
rect 16448 36116 16454 36168
rect 16482 36116 16488 36168
rect 16540 36156 16546 36168
rect 17129 36159 17187 36165
rect 16540 36128 16585 36156
rect 16540 36116 16546 36128
rect 17129 36125 17141 36159
rect 17175 36125 17187 36159
rect 17770 36156 17776 36168
rect 17731 36128 17776 36156
rect 17129 36119 17187 36125
rect 3016 36060 3280 36088
rect 3016 36048 3022 36060
rect 4614 36048 4620 36100
rect 4672 36088 4678 36100
rect 5629 36091 5687 36097
rect 5629 36088 5641 36091
rect 4672 36060 5641 36088
rect 4672 36048 4678 36060
rect 5629 36057 5641 36060
rect 5675 36057 5687 36091
rect 5629 36051 5687 36057
rect 5810 36048 5816 36100
rect 5868 36088 5874 36100
rect 7101 36091 7159 36097
rect 7101 36088 7113 36091
rect 5868 36060 7113 36088
rect 5868 36048 5874 36060
rect 7101 36057 7113 36060
rect 7147 36088 7159 36091
rect 9766 36088 9772 36100
rect 7147 36060 9772 36088
rect 7147 36057 7159 36060
rect 7101 36051 7159 36057
rect 9766 36048 9772 36060
rect 9824 36048 9830 36100
rect 9950 36088 9956 36100
rect 9911 36060 9956 36088
rect 9950 36048 9956 36060
rect 10008 36048 10014 36100
rect 12253 36091 12311 36097
rect 12253 36057 12265 36091
rect 12299 36088 12311 36091
rect 12526 36088 12532 36100
rect 12299 36060 12532 36088
rect 12299 36057 12311 36060
rect 12253 36051 12311 36057
rect 12526 36048 12532 36060
rect 12584 36048 12590 36100
rect 13173 36091 13231 36097
rect 13173 36057 13185 36091
rect 13219 36088 13231 36091
rect 13354 36088 13360 36100
rect 13219 36060 13360 36088
rect 13219 36057 13231 36060
rect 13173 36051 13231 36057
rect 13354 36048 13360 36060
rect 13412 36048 13418 36100
rect 14182 36048 14188 36100
rect 14240 36088 14246 36100
rect 15562 36088 15568 36100
rect 14240 36060 14398 36088
rect 15523 36060 15568 36088
rect 14240 36048 14246 36060
rect 15562 36048 15568 36060
rect 15620 36048 15626 36100
rect 9858 35980 9864 36032
rect 9916 36020 9922 36032
rect 10686 36020 10692 36032
rect 9916 35992 10692 36020
rect 9916 35980 9922 35992
rect 10686 35980 10692 35992
rect 10744 35980 10750 36032
rect 12434 35980 12440 36032
rect 12492 36020 12498 36032
rect 12805 36023 12863 36029
rect 12805 36020 12817 36023
rect 12492 35992 12817 36020
rect 12492 35980 12498 35992
rect 12805 35989 12817 35992
rect 12851 35989 12863 36023
rect 14090 36020 14096 36032
rect 14051 35992 14096 36020
rect 12805 35983 12863 35989
rect 14090 35980 14096 35992
rect 14148 35980 14154 36032
rect 15654 35980 15660 36032
rect 15712 36020 15718 36032
rect 16301 36023 16359 36029
rect 16301 36020 16313 36023
rect 15712 35992 16313 36020
rect 15712 35980 15718 35992
rect 16301 35989 16313 35992
rect 16347 35989 16359 36023
rect 17144 36020 17172 36119
rect 17770 36116 17776 36128
rect 17828 36116 17834 36168
rect 18506 36156 18512 36168
rect 18467 36128 18512 36156
rect 18506 36116 18512 36128
rect 18564 36116 18570 36168
rect 21174 36116 21180 36168
rect 21232 36156 21238 36168
rect 21545 36159 21603 36165
rect 21545 36156 21557 36159
rect 21232 36128 21557 36156
rect 21232 36116 21238 36128
rect 21545 36125 21557 36128
rect 21591 36125 21603 36159
rect 21545 36119 21603 36125
rect 22646 36116 22652 36168
rect 22704 36156 22710 36168
rect 23017 36159 23075 36165
rect 23017 36156 23029 36159
rect 22704 36128 23029 36156
rect 22704 36116 22710 36128
rect 23017 36125 23029 36128
rect 23063 36125 23075 36159
rect 24578 36156 24584 36168
rect 24539 36128 24584 36156
rect 23017 36119 23075 36125
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 25225 36159 25283 36165
rect 25225 36125 25237 36159
rect 25271 36156 25283 36159
rect 25314 36156 25320 36168
rect 25271 36128 25320 36156
rect 25271 36125 25283 36128
rect 25225 36119 25283 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 28445 36159 28503 36165
rect 28445 36125 28457 36159
rect 28491 36125 28503 36159
rect 28445 36119 28503 36125
rect 18601 36091 18659 36097
rect 18601 36057 18613 36091
rect 18647 36088 18659 36091
rect 19429 36091 19487 36097
rect 19429 36088 19441 36091
rect 18647 36060 19441 36088
rect 18647 36057 18659 36060
rect 18601 36051 18659 36057
rect 19429 36057 19441 36060
rect 19475 36057 19487 36091
rect 22370 36088 22376 36100
rect 22331 36060 22376 36088
rect 19429 36051 19487 36057
rect 22370 36048 22376 36060
rect 22428 36048 22434 36100
rect 28460 36088 28488 36119
rect 28534 36116 28540 36168
rect 28592 36156 28598 36168
rect 28629 36159 28687 36165
rect 28629 36156 28641 36159
rect 28592 36128 28641 36156
rect 28592 36116 28598 36128
rect 28629 36125 28641 36128
rect 28675 36125 28687 36159
rect 28629 36119 28687 36125
rect 28994 36116 29000 36168
rect 29052 36156 29058 36168
rect 29549 36159 29607 36165
rect 29549 36156 29561 36159
rect 29052 36128 29561 36156
rect 29052 36116 29058 36128
rect 29549 36125 29561 36128
rect 29595 36125 29607 36159
rect 29549 36119 29607 36125
rect 34149 36159 34207 36165
rect 34149 36125 34161 36159
rect 34195 36156 34207 36159
rect 34606 36156 34612 36168
rect 34195 36128 34612 36156
rect 34195 36125 34207 36128
rect 34149 36119 34207 36125
rect 34606 36116 34612 36128
rect 34664 36116 34670 36168
rect 34698 36116 34704 36168
rect 34756 36156 34762 36168
rect 35805 36159 35863 36165
rect 34756 36128 34801 36156
rect 34756 36116 34762 36128
rect 35805 36125 35817 36159
rect 35851 36156 35863 36159
rect 36265 36159 36323 36165
rect 36265 36156 36277 36159
rect 35851 36128 36277 36156
rect 35851 36125 35863 36128
rect 35805 36119 35863 36125
rect 36265 36125 36277 36128
rect 36311 36125 36323 36159
rect 36265 36119 36323 36125
rect 28810 36088 28816 36100
rect 28460 36060 28816 36088
rect 28810 36048 28816 36060
rect 28868 36048 28874 36100
rect 31846 36088 31852 36100
rect 31807 36060 31852 36088
rect 31846 36048 31852 36060
rect 31904 36048 31910 36100
rect 36449 36091 36507 36097
rect 36449 36057 36461 36091
rect 36495 36088 36507 36091
rect 37458 36088 37464 36100
rect 36495 36060 37464 36088
rect 36495 36057 36507 36060
rect 36449 36051 36507 36057
rect 37458 36048 37464 36060
rect 37516 36048 37522 36100
rect 20898 36020 20904 36032
rect 17144 35992 20904 36020
rect 16301 35983 16359 35989
rect 20898 35980 20904 35992
rect 20956 35980 20962 36032
rect 25038 35980 25044 36032
rect 25096 36020 25102 36032
rect 25133 36023 25191 36029
rect 25133 36020 25145 36023
rect 25096 35992 25145 36020
rect 25096 35980 25102 35992
rect 25133 35989 25145 35992
rect 25179 35989 25191 36023
rect 25133 35983 25191 35989
rect 28442 35980 28448 36032
rect 28500 36020 28506 36032
rect 28537 36023 28595 36029
rect 28537 36020 28549 36023
rect 28500 35992 28549 36020
rect 28500 35980 28506 35992
rect 28537 35989 28549 35992
rect 28583 35989 28595 36023
rect 28537 35983 28595 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 4525 35819 4583 35825
rect 4525 35785 4537 35819
rect 4571 35816 4583 35819
rect 5534 35816 5540 35828
rect 4571 35788 5540 35816
rect 4571 35785 4583 35788
rect 4525 35779 4583 35785
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 9122 35776 9128 35828
rect 9180 35816 9186 35828
rect 9674 35816 9680 35828
rect 9180 35788 9680 35816
rect 9180 35776 9186 35788
rect 9674 35776 9680 35788
rect 9732 35776 9738 35828
rect 9769 35819 9827 35825
rect 9769 35785 9781 35819
rect 9815 35816 9827 35819
rect 9950 35816 9956 35828
rect 9815 35788 9956 35816
rect 9815 35785 9827 35788
rect 9769 35779 9827 35785
rect 9950 35776 9956 35788
rect 10008 35776 10014 35828
rect 10413 35819 10471 35825
rect 10413 35785 10425 35819
rect 10459 35816 10471 35819
rect 11698 35816 11704 35828
rect 10459 35788 11704 35816
rect 10459 35785 10471 35788
rect 10413 35779 10471 35785
rect 11698 35776 11704 35788
rect 11756 35776 11762 35828
rect 14829 35819 14887 35825
rect 14829 35785 14841 35819
rect 14875 35816 14887 35819
rect 15562 35816 15568 35828
rect 14875 35788 15568 35816
rect 14875 35785 14887 35788
rect 14829 35779 14887 35785
rect 15562 35776 15568 35788
rect 15620 35776 15626 35828
rect 21726 35776 21732 35828
rect 21784 35816 21790 35828
rect 21913 35819 21971 35825
rect 21913 35816 21925 35819
rect 21784 35788 21925 35816
rect 21784 35776 21790 35788
rect 21913 35785 21925 35788
rect 21959 35785 21971 35819
rect 21913 35779 21971 35785
rect 27157 35819 27215 35825
rect 27157 35785 27169 35819
rect 27203 35816 27215 35819
rect 27246 35816 27252 35828
rect 27203 35788 27252 35816
rect 27203 35785 27215 35788
rect 27157 35779 27215 35785
rect 27246 35776 27252 35788
rect 27304 35776 27310 35828
rect 29546 35776 29552 35828
rect 29604 35816 29610 35828
rect 30193 35819 30251 35825
rect 30193 35816 30205 35819
rect 29604 35788 30205 35816
rect 29604 35776 29610 35788
rect 30193 35785 30205 35788
rect 30239 35785 30251 35819
rect 30193 35779 30251 35785
rect 31846 35776 31852 35828
rect 31904 35816 31910 35828
rect 32217 35819 32275 35825
rect 32217 35816 32229 35819
rect 31904 35788 32229 35816
rect 31904 35776 31910 35788
rect 32217 35785 32229 35788
rect 32263 35785 32275 35819
rect 32217 35779 32275 35785
rect 32582 35776 32588 35828
rect 32640 35816 32646 35828
rect 32861 35819 32919 35825
rect 32861 35816 32873 35819
rect 32640 35788 32873 35816
rect 32640 35776 32646 35788
rect 32861 35785 32873 35788
rect 32907 35785 32919 35819
rect 37458 35816 37464 35828
rect 37419 35788 37464 35816
rect 32861 35779 32919 35785
rect 37458 35776 37464 35788
rect 37516 35776 37522 35828
rect 5353 35751 5411 35757
rect 5353 35717 5365 35751
rect 5399 35748 5411 35751
rect 7282 35748 7288 35760
rect 5399 35720 7288 35748
rect 5399 35717 5411 35720
rect 5353 35711 5411 35717
rect 7282 35708 7288 35720
rect 7340 35708 7346 35760
rect 12526 35708 12532 35760
rect 12584 35708 12590 35760
rect 14553 35751 14611 35757
rect 14553 35717 14565 35751
rect 14599 35748 14611 35751
rect 16025 35751 16083 35757
rect 16025 35748 16037 35751
rect 14599 35720 16037 35748
rect 14599 35717 14611 35720
rect 14553 35711 14611 35717
rect 16025 35717 16037 35720
rect 16071 35717 16083 35751
rect 16025 35711 16083 35717
rect 21358 35708 21364 35760
rect 21416 35748 21422 35760
rect 35069 35751 35127 35757
rect 21416 35720 32628 35748
rect 21416 35708 21422 35720
rect 32600 35692 32628 35720
rect 35069 35717 35081 35751
rect 35115 35748 35127 35751
rect 35894 35748 35900 35760
rect 35115 35720 35900 35748
rect 35115 35717 35127 35720
rect 35069 35711 35127 35717
rect 35894 35708 35900 35720
rect 35952 35708 35958 35760
rect 36725 35751 36783 35757
rect 36725 35717 36737 35751
rect 36771 35748 36783 35751
rect 38010 35748 38016 35760
rect 36771 35720 38016 35748
rect 36771 35717 36783 35720
rect 36725 35711 36783 35717
rect 38010 35708 38016 35720
rect 38068 35708 38074 35760
rect 4617 35683 4675 35689
rect 4617 35649 4629 35683
rect 4663 35649 4675 35683
rect 4617 35643 4675 35649
rect 5721 35683 5779 35689
rect 5721 35649 5733 35683
rect 5767 35680 5779 35683
rect 6454 35680 6460 35692
rect 5767 35652 6460 35680
rect 5767 35649 5779 35652
rect 5721 35643 5779 35649
rect 1762 35612 1768 35624
rect 1723 35584 1768 35612
rect 1762 35572 1768 35584
rect 1820 35572 1826 35624
rect 1949 35615 2007 35621
rect 1949 35581 1961 35615
rect 1995 35612 2007 35615
rect 2222 35612 2228 35624
rect 1995 35584 2228 35612
rect 1995 35581 2007 35584
rect 1949 35575 2007 35581
rect 2222 35572 2228 35584
rect 2280 35572 2286 35624
rect 2774 35612 2780 35624
rect 2735 35584 2780 35612
rect 2774 35572 2780 35584
rect 2832 35572 2838 35624
rect 4632 35612 4660 35643
rect 6454 35640 6460 35652
rect 6512 35640 6518 35692
rect 8386 35680 8392 35692
rect 8347 35652 8392 35680
rect 8386 35640 8392 35652
rect 8444 35640 8450 35692
rect 9677 35683 9735 35689
rect 9677 35649 9689 35683
rect 9723 35680 9735 35683
rect 9858 35680 9864 35692
rect 9723 35652 9864 35680
rect 9723 35649 9735 35652
rect 9677 35643 9735 35649
rect 9858 35640 9864 35652
rect 9916 35640 9922 35692
rect 10502 35680 10508 35692
rect 10463 35652 10508 35680
rect 10502 35640 10508 35652
rect 10560 35640 10566 35692
rect 14090 35640 14096 35692
rect 14148 35680 14154 35692
rect 14366 35689 14372 35692
rect 14185 35683 14243 35689
rect 14185 35680 14197 35683
rect 14148 35652 14197 35680
rect 14148 35640 14154 35652
rect 14185 35649 14197 35652
rect 14231 35649 14243 35683
rect 14185 35643 14243 35649
rect 14343 35683 14372 35689
rect 14343 35649 14355 35683
rect 14343 35643 14372 35649
rect 14366 35640 14372 35643
rect 14424 35640 14430 35692
rect 14458 35640 14464 35692
rect 14516 35680 14522 35692
rect 14645 35683 14703 35689
rect 14516 35652 14561 35680
rect 14516 35640 14522 35652
rect 14645 35649 14657 35683
rect 14691 35680 14703 35683
rect 15102 35680 15108 35692
rect 14691 35652 15108 35680
rect 14691 35649 14703 35652
rect 14645 35643 14703 35649
rect 15102 35640 15108 35652
rect 15160 35640 15166 35692
rect 15286 35680 15292 35692
rect 15247 35652 15292 35680
rect 15286 35640 15292 35652
rect 15344 35640 15350 35692
rect 15473 35683 15531 35689
rect 15473 35649 15485 35683
rect 15519 35649 15531 35683
rect 15930 35680 15936 35692
rect 15891 35652 15936 35680
rect 15473 35643 15531 35649
rect 5994 35612 6000 35624
rect 4632 35584 6000 35612
rect 5994 35572 6000 35584
rect 6052 35572 6058 35624
rect 7190 35612 7196 35624
rect 7151 35584 7196 35612
rect 7190 35572 7196 35584
rect 7248 35572 7254 35624
rect 11514 35572 11520 35624
rect 11572 35612 11578 35624
rect 11701 35615 11759 35621
rect 11701 35612 11713 35615
rect 11572 35584 11713 35612
rect 11572 35572 11578 35584
rect 11701 35581 11713 35584
rect 11747 35581 11759 35615
rect 11974 35612 11980 35624
rect 11935 35584 11980 35612
rect 11701 35575 11759 35581
rect 11974 35572 11980 35584
rect 12032 35572 12038 35624
rect 13814 35572 13820 35624
rect 13872 35612 13878 35624
rect 15488 35612 15516 35643
rect 15930 35640 15936 35652
rect 15988 35640 15994 35692
rect 16390 35640 16396 35692
rect 16448 35680 16454 35692
rect 17037 35683 17095 35689
rect 17037 35680 17049 35683
rect 16448 35652 17049 35680
rect 16448 35640 16454 35652
rect 17037 35649 17049 35652
rect 17083 35649 17095 35683
rect 19334 35680 19340 35692
rect 18446 35652 19340 35680
rect 17037 35643 17095 35649
rect 19334 35640 19340 35652
rect 19392 35640 19398 35692
rect 19518 35680 19524 35692
rect 19479 35652 19524 35680
rect 19518 35640 19524 35652
rect 19576 35680 19582 35692
rect 20254 35680 20260 35692
rect 19576 35652 20260 35680
rect 19576 35640 19582 35652
rect 20254 35640 20260 35652
rect 20312 35640 20318 35692
rect 20441 35683 20499 35689
rect 20441 35649 20453 35683
rect 20487 35680 20499 35683
rect 20714 35680 20720 35692
rect 20487 35652 20720 35680
rect 20487 35649 20499 35652
rect 20441 35643 20499 35649
rect 13872 35584 15516 35612
rect 17313 35615 17371 35621
rect 13872 35572 13878 35584
rect 17313 35581 17325 35615
rect 17359 35612 17371 35615
rect 17678 35612 17684 35624
rect 17359 35584 17684 35612
rect 17359 35581 17371 35584
rect 17313 35575 17371 35581
rect 17678 35572 17684 35584
rect 17736 35572 17742 35624
rect 15289 35547 15347 35553
rect 15289 35544 15301 35547
rect 13372 35516 15301 35544
rect 11238 35436 11244 35488
rect 11296 35476 11302 35488
rect 13372 35476 13400 35516
rect 15289 35513 15301 35516
rect 15335 35513 15347 35547
rect 15289 35507 15347 35513
rect 19705 35547 19763 35553
rect 19705 35513 19717 35547
rect 19751 35544 19763 35547
rect 20456 35544 20484 35643
rect 20714 35640 20720 35652
rect 20772 35680 20778 35692
rect 21174 35680 21180 35692
rect 20772 35652 21180 35680
rect 20772 35640 20778 35652
rect 21174 35640 21180 35652
rect 21232 35640 21238 35692
rect 22002 35680 22008 35692
rect 21963 35652 22008 35680
rect 22002 35640 22008 35652
rect 22060 35640 22066 35692
rect 22646 35680 22652 35692
rect 22607 35652 22652 35680
rect 22646 35640 22652 35652
rect 22704 35640 22710 35692
rect 25317 35683 25375 35689
rect 25317 35649 25329 35683
rect 25363 35680 25375 35683
rect 25498 35680 25504 35692
rect 25363 35652 25504 35680
rect 25363 35649 25375 35652
rect 25317 35643 25375 35649
rect 25498 35640 25504 35652
rect 25556 35640 25562 35692
rect 26145 35683 26203 35689
rect 26145 35649 26157 35683
rect 26191 35680 26203 35683
rect 26970 35680 26976 35692
rect 26191 35652 26976 35680
rect 26191 35649 26203 35652
rect 26145 35643 26203 35649
rect 26970 35640 26976 35652
rect 27028 35640 27034 35692
rect 27338 35680 27344 35692
rect 27299 35652 27344 35680
rect 27338 35640 27344 35652
rect 27396 35640 27402 35692
rect 27798 35680 27804 35692
rect 27759 35652 27804 35680
rect 27798 35640 27804 35652
rect 27856 35640 27862 35692
rect 30098 35680 30104 35692
rect 30059 35652 30104 35680
rect 30098 35640 30104 35652
rect 30156 35640 30162 35692
rect 32214 35640 32220 35692
rect 32272 35680 32278 35692
rect 32309 35683 32367 35689
rect 32309 35680 32321 35683
rect 32272 35652 32321 35680
rect 32272 35640 32278 35652
rect 32309 35649 32321 35652
rect 32355 35649 32367 35683
rect 32309 35643 32367 35649
rect 32582 35640 32588 35692
rect 32640 35680 32646 35692
rect 32953 35683 33011 35689
rect 32953 35680 32965 35683
rect 32640 35652 32965 35680
rect 32640 35640 32646 35652
rect 32953 35649 32965 35652
rect 32999 35649 33011 35683
rect 32953 35643 33011 35649
rect 34606 35640 34612 35692
rect 34664 35680 34670 35692
rect 34885 35683 34943 35689
rect 34885 35680 34897 35683
rect 34664 35652 34897 35680
rect 34664 35640 34670 35652
rect 34885 35649 34897 35652
rect 34931 35649 34943 35683
rect 34885 35643 34943 35649
rect 37369 35683 37427 35689
rect 37369 35649 37381 35683
rect 37415 35680 37427 35683
rect 38378 35680 38384 35692
rect 37415 35652 38384 35680
rect 37415 35649 37427 35652
rect 37369 35643 37427 35649
rect 20806 35612 20812 35624
rect 20767 35584 20812 35612
rect 20806 35572 20812 35584
rect 20864 35572 20870 35624
rect 22830 35612 22836 35624
rect 22791 35584 22836 35612
rect 22830 35572 22836 35584
rect 22888 35572 22894 35624
rect 23198 35612 23204 35624
rect 23159 35584 23204 35612
rect 23198 35572 23204 35584
rect 23256 35572 23262 35624
rect 27982 35612 27988 35624
rect 27943 35584 27988 35612
rect 27982 35572 27988 35584
rect 28040 35572 28046 35624
rect 28350 35612 28356 35624
rect 28311 35584 28356 35612
rect 28350 35572 28356 35584
rect 28408 35572 28414 35624
rect 19751 35516 20484 35544
rect 19751 35513 19763 35516
rect 19705 35507 19763 35513
rect 20990 35504 20996 35556
rect 21048 35544 21054 35556
rect 21818 35544 21824 35556
rect 21048 35516 21824 35544
rect 21048 35504 21054 35516
rect 21818 35504 21824 35516
rect 21876 35544 21882 35556
rect 37384 35544 37412 35643
rect 38378 35640 38384 35652
rect 38436 35640 38442 35692
rect 21876 35516 37412 35544
rect 21876 35504 21882 35516
rect 11296 35448 13400 35476
rect 13449 35479 13507 35485
rect 11296 35436 11302 35448
rect 13449 35445 13461 35479
rect 13495 35476 13507 35479
rect 13538 35476 13544 35488
rect 13495 35448 13544 35476
rect 13495 35445 13507 35448
rect 13449 35439 13507 35445
rect 13538 35436 13544 35448
rect 13596 35436 13602 35488
rect 13630 35436 13636 35488
rect 13688 35476 13694 35488
rect 14366 35476 14372 35488
rect 13688 35448 14372 35476
rect 13688 35436 13694 35448
rect 14366 35436 14372 35448
rect 14424 35476 14430 35488
rect 17034 35476 17040 35488
rect 14424 35448 17040 35476
rect 14424 35436 14430 35448
rect 17034 35436 17040 35448
rect 17092 35436 17098 35488
rect 18322 35436 18328 35488
rect 18380 35476 18386 35488
rect 18785 35479 18843 35485
rect 18785 35476 18797 35479
rect 18380 35448 18797 35476
rect 18380 35436 18386 35448
rect 18785 35445 18797 35448
rect 18831 35445 18843 35479
rect 25130 35476 25136 35488
rect 25091 35448 25136 35476
rect 18785 35439 18843 35445
rect 25130 35436 25136 35448
rect 25188 35436 25194 35488
rect 26053 35479 26111 35485
rect 26053 35445 26065 35479
rect 26099 35476 26111 35479
rect 26234 35476 26240 35488
rect 26099 35448 26240 35476
rect 26099 35445 26111 35448
rect 26053 35439 26111 35445
rect 26234 35436 26240 35448
rect 26292 35436 26298 35488
rect 26878 35436 26884 35488
rect 26936 35476 26942 35488
rect 36722 35476 36728 35488
rect 26936 35448 36728 35476
rect 26936 35436 26942 35448
rect 36722 35436 36728 35448
rect 36780 35436 36786 35488
rect 36814 35436 36820 35488
rect 36872 35476 36878 35488
rect 38010 35476 38016 35488
rect 36872 35448 38016 35476
rect 36872 35436 36878 35448
rect 38010 35436 38016 35448
rect 38068 35436 38074 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 4065 35275 4123 35281
rect 4065 35241 4077 35275
rect 4111 35272 4123 35275
rect 4614 35272 4620 35284
rect 4111 35244 4620 35272
rect 4111 35241 4123 35244
rect 4065 35235 4123 35241
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 11974 35232 11980 35284
rect 12032 35272 12038 35284
rect 12253 35275 12311 35281
rect 12253 35272 12265 35275
rect 12032 35244 12265 35272
rect 12032 35232 12038 35244
rect 12253 35241 12265 35244
rect 12299 35241 12311 35275
rect 12253 35235 12311 35241
rect 12526 35232 12532 35284
rect 12584 35272 12590 35284
rect 13449 35275 13507 35281
rect 13449 35272 13461 35275
rect 12584 35244 13461 35272
rect 12584 35232 12590 35244
rect 13449 35241 13461 35244
rect 13495 35272 13507 35275
rect 15286 35272 15292 35284
rect 13495 35244 15292 35272
rect 13495 35241 13507 35244
rect 13449 35235 13507 35241
rect 15286 35232 15292 35244
rect 15344 35232 15350 35284
rect 17678 35272 17684 35284
rect 17639 35244 17684 35272
rect 17678 35232 17684 35244
rect 17736 35232 17742 35284
rect 19334 35272 19340 35284
rect 19295 35244 19340 35272
rect 19334 35232 19340 35244
rect 19392 35232 19398 35284
rect 24578 35232 24584 35284
rect 24636 35272 24642 35284
rect 27338 35272 27344 35284
rect 24636 35244 26740 35272
rect 27299 35244 27344 35272
rect 24636 35232 24642 35244
rect 14458 35204 14464 35216
rect 12636 35176 14464 35204
rect 2685 35139 2743 35145
rect 2685 35105 2697 35139
rect 2731 35136 2743 35139
rect 2866 35136 2872 35148
rect 2731 35108 2872 35136
rect 2731 35105 2743 35108
rect 2685 35099 2743 35105
rect 2866 35096 2872 35108
rect 2924 35096 2930 35148
rect 10686 35096 10692 35148
rect 10744 35136 10750 35148
rect 10744 35108 11560 35136
rect 10744 35096 10750 35108
rect 3234 35028 3240 35080
rect 3292 35068 3298 35080
rect 3973 35071 4031 35077
rect 3292 35040 3337 35068
rect 3292 35028 3298 35040
rect 3973 35037 3985 35071
rect 4019 35068 4031 35071
rect 5810 35068 5816 35080
rect 4019 35040 5488 35068
rect 5771 35040 5816 35068
rect 4019 35037 4031 35040
rect 3973 35031 4031 35037
rect 5460 35012 5488 35040
rect 5810 35028 5816 35040
rect 5868 35028 5874 35080
rect 6454 35068 6460 35080
rect 6415 35040 6460 35068
rect 6454 35028 6460 35040
rect 6512 35028 6518 35080
rect 8478 35028 8484 35080
rect 8536 35068 8542 35080
rect 8941 35071 8999 35077
rect 8941 35068 8953 35071
rect 8536 35040 8953 35068
rect 8536 35028 8542 35040
rect 8941 35037 8953 35040
rect 8987 35037 8999 35071
rect 11238 35068 11244 35080
rect 11199 35040 11244 35068
rect 8941 35031 8999 35037
rect 11238 35028 11244 35040
rect 11296 35028 11302 35080
rect 11532 35077 11560 35108
rect 11517 35071 11575 35077
rect 11517 35037 11529 35071
rect 11563 35068 11575 35071
rect 12158 35068 12164 35080
rect 11563 35040 12164 35068
rect 11563 35037 11575 35040
rect 11517 35031 11575 35037
rect 12158 35028 12164 35040
rect 12216 35028 12222 35080
rect 12434 35028 12440 35080
rect 12492 35068 12498 35080
rect 12492 35040 12537 35068
rect 12492 35028 12498 35040
rect 2866 34960 2872 35012
rect 2924 35000 2930 35012
rect 3053 35003 3111 35009
rect 3053 35000 3065 35003
rect 2924 34972 3065 35000
rect 2924 34960 2930 34972
rect 3053 34969 3065 34972
rect 3099 34969 3111 35003
rect 5442 35000 5448 35012
rect 5403 34972 5448 35000
rect 3053 34963 3111 34969
rect 5442 34960 5448 34972
rect 5500 34960 5506 35012
rect 6178 34960 6184 35012
rect 6236 35000 6242 35012
rect 6825 35003 6883 35009
rect 6825 35000 6837 35003
rect 6236 34972 6837 35000
rect 6236 34960 6242 34972
rect 6825 34969 6837 34972
rect 6871 35000 6883 35003
rect 8846 35000 8852 35012
rect 6871 34972 8852 35000
rect 6871 34969 6883 34972
rect 6825 34963 6883 34969
rect 8846 34960 8852 34972
rect 8904 34960 8910 35012
rect 9217 35003 9275 35009
rect 9217 34969 9229 35003
rect 9263 34969 9275 35003
rect 10778 35000 10784 35012
rect 10442 34972 10784 35000
rect 9217 34963 9275 34969
rect 9232 34932 9260 34963
rect 10778 34960 10784 34972
rect 10836 34960 10842 35012
rect 11333 35003 11391 35009
rect 11333 34969 11345 35003
rect 11379 35000 11391 35003
rect 11974 35000 11980 35012
rect 11379 34972 11980 35000
rect 11379 34969 11391 34972
rect 11333 34963 11391 34969
rect 11974 34960 11980 34972
rect 12032 34960 12038 35012
rect 12526 35000 12532 35012
rect 12487 34972 12532 35000
rect 12526 34960 12532 34972
rect 12584 34960 12590 35012
rect 12636 35009 12664 35176
rect 14458 35164 14464 35176
rect 14516 35204 14522 35216
rect 16206 35204 16212 35216
rect 14516 35176 16212 35204
rect 14516 35164 14522 35176
rect 16206 35164 16212 35176
rect 16264 35164 16270 35216
rect 18138 35204 18144 35216
rect 16408 35176 18144 35204
rect 12897 35139 12955 35145
rect 12897 35105 12909 35139
rect 12943 35136 12955 35139
rect 12943 35108 13584 35136
rect 12943 35105 12955 35108
rect 12897 35099 12955 35105
rect 13556 35080 13584 35108
rect 14090 35096 14096 35148
rect 14148 35136 14154 35148
rect 15105 35139 15163 35145
rect 15105 35136 15117 35139
rect 14148 35108 15117 35136
rect 14148 35096 14154 35108
rect 15105 35105 15117 35108
rect 15151 35105 15163 35139
rect 15657 35139 15715 35145
rect 15657 35136 15669 35139
rect 15105 35099 15163 35105
rect 15212 35108 15669 35136
rect 13354 35068 13360 35080
rect 13315 35040 13360 35068
rect 13354 35028 13360 35040
rect 13412 35028 13418 35080
rect 13538 35068 13544 35080
rect 13499 35040 13544 35068
rect 13538 35028 13544 35040
rect 13596 35028 13602 35080
rect 13906 35028 13912 35080
rect 13964 35068 13970 35080
rect 14277 35071 14335 35077
rect 14277 35068 14289 35071
rect 13964 35040 14289 35068
rect 13964 35028 13970 35040
rect 14277 35037 14289 35040
rect 14323 35037 14335 35071
rect 14277 35031 14335 35037
rect 12621 35003 12679 35009
rect 12621 34969 12633 35003
rect 12667 34969 12679 35003
rect 12621 34963 12679 34969
rect 10594 34932 10600 34944
rect 9232 34904 10600 34932
rect 10594 34892 10600 34904
rect 10652 34892 10658 34944
rect 10686 34892 10692 34944
rect 10744 34932 10750 34944
rect 11698 34932 11704 34944
rect 10744 34904 10789 34932
rect 11659 34904 11704 34932
rect 10744 34892 10750 34904
rect 11698 34892 11704 34904
rect 11756 34892 11762 34944
rect 11882 34892 11888 34944
rect 11940 34932 11946 34944
rect 12636 34932 12664 34963
rect 12710 34960 12716 35012
rect 12768 35009 12774 35012
rect 12768 35003 12817 35009
rect 12768 34969 12771 35003
rect 12805 35000 12817 35003
rect 13372 35000 13400 35028
rect 14458 35000 14464 35012
rect 12805 34972 13308 35000
rect 13372 34972 14464 35000
rect 12805 34969 12817 34972
rect 12768 34963 12817 34969
rect 12768 34960 12774 34963
rect 11940 34904 12664 34932
rect 13280 34932 13308 34972
rect 14458 34960 14464 34972
rect 14516 35000 14522 35012
rect 15212 35000 15240 35108
rect 15657 35105 15669 35108
rect 15703 35136 15715 35139
rect 15930 35136 15936 35148
rect 15703 35108 15936 35136
rect 15703 35105 15715 35108
rect 15657 35099 15715 35105
rect 15930 35096 15936 35108
rect 15988 35096 15994 35148
rect 15286 35028 15292 35080
rect 15344 35068 15350 35080
rect 15473 35071 15531 35077
rect 15473 35068 15485 35071
rect 15344 35040 15485 35068
rect 15344 35028 15350 35040
rect 15473 35037 15485 35040
rect 15519 35068 15531 35071
rect 16298 35068 16304 35080
rect 15519 35040 16304 35068
rect 15519 35037 15531 35040
rect 15473 35031 15531 35037
rect 16298 35028 16304 35040
rect 16356 35068 16362 35080
rect 16408 35077 16436 35176
rect 18138 35164 18144 35176
rect 18196 35164 18202 35216
rect 17037 35139 17095 35145
rect 17037 35105 17049 35139
rect 17083 35136 17095 35139
rect 18322 35136 18328 35148
rect 17083 35108 18328 35136
rect 17083 35105 17095 35108
rect 17037 35099 17095 35105
rect 16393 35071 16451 35077
rect 16393 35068 16405 35071
rect 16356 35040 16405 35068
rect 16356 35028 16362 35040
rect 16393 35037 16405 35040
rect 16439 35037 16451 35071
rect 16393 35031 16451 35037
rect 16577 35071 16635 35077
rect 16577 35037 16589 35071
rect 16623 35068 16635 35071
rect 17052 35068 17080 35099
rect 18322 35096 18328 35108
rect 18380 35096 18386 35148
rect 24854 35136 24860 35148
rect 24767 35108 24860 35136
rect 24854 35096 24860 35108
rect 24912 35136 24918 35148
rect 26142 35136 26148 35148
rect 24912 35108 26148 35136
rect 24912 35096 24918 35108
rect 26142 35096 26148 35108
rect 26200 35096 26206 35148
rect 16623 35040 17080 35068
rect 17497 35071 17555 35077
rect 16623 35037 16635 35040
rect 16577 35031 16635 35037
rect 17497 35037 17509 35071
rect 17543 35068 17555 35071
rect 18509 35071 18567 35077
rect 18509 35068 18521 35071
rect 17543 35040 18521 35068
rect 17543 35037 17555 35040
rect 17497 35031 17555 35037
rect 18509 35037 18521 35040
rect 18555 35037 18567 35071
rect 19426 35068 19432 35080
rect 19339 35040 19432 35068
rect 18509 35031 18567 35037
rect 14516 34972 15240 35000
rect 14516 34960 14522 34972
rect 15378 34960 15384 35012
rect 15436 35000 15442 35012
rect 16592 35000 16620 35031
rect 19426 35028 19432 35040
rect 19484 35068 19490 35080
rect 20162 35068 20168 35080
rect 19484 35040 20168 35068
rect 19484 35028 19490 35040
rect 20162 35028 20168 35040
rect 20220 35028 20226 35080
rect 20714 35068 20720 35080
rect 20675 35040 20720 35068
rect 20714 35028 20720 35040
rect 20772 35028 20778 35080
rect 23845 35071 23903 35077
rect 23845 35037 23857 35071
rect 23891 35037 23903 35071
rect 23845 35031 23903 35037
rect 15436 34972 16620 35000
rect 15436 34960 15442 34972
rect 17034 34960 17040 35012
rect 17092 35000 17098 35012
rect 17175 35003 17233 35009
rect 17175 35000 17187 35003
rect 17092 34972 17187 35000
rect 17092 34960 17098 34972
rect 17175 34969 17187 34972
rect 17221 34969 17233 35003
rect 17175 34963 17233 34969
rect 17313 35003 17371 35009
rect 17313 34969 17325 35003
rect 17359 34969 17371 35003
rect 17313 34963 17371 34969
rect 13630 34932 13636 34944
rect 13280 34904 13636 34932
rect 11940 34892 11946 34904
rect 13630 34892 13636 34904
rect 13688 34892 13694 34944
rect 13814 34892 13820 34944
rect 13872 34932 13878 34944
rect 14185 34935 14243 34941
rect 14185 34932 14197 34935
rect 13872 34904 14197 34932
rect 13872 34892 13878 34904
rect 14185 34901 14197 34904
rect 14231 34901 14243 34935
rect 14185 34895 14243 34901
rect 15194 34892 15200 34944
rect 15252 34932 15258 34944
rect 15289 34935 15347 34941
rect 15289 34932 15301 34935
rect 15252 34904 15301 34932
rect 15252 34892 15258 34904
rect 15289 34901 15301 34904
rect 15335 34932 15347 34935
rect 15470 34932 15476 34944
rect 15335 34904 15476 34932
rect 15335 34901 15347 34904
rect 15289 34895 15347 34901
rect 15470 34892 15476 34904
rect 15528 34892 15534 34944
rect 16577 34935 16635 34941
rect 16577 34901 16589 34935
rect 16623 34932 16635 34935
rect 16850 34932 16856 34944
rect 16623 34904 16856 34932
rect 16623 34901 16635 34904
rect 16577 34895 16635 34901
rect 16850 34892 16856 34904
rect 16908 34932 16914 34944
rect 17328 34932 17356 34963
rect 17402 34960 17408 35012
rect 17460 35000 17466 35012
rect 18138 35000 18144 35012
rect 17460 34972 17505 35000
rect 18099 34972 18144 35000
rect 17460 34960 17466 34972
rect 18138 34960 18144 34972
rect 18196 34960 18202 35012
rect 18322 35000 18328 35012
rect 18283 34972 18328 35000
rect 18322 34960 18328 34972
rect 18380 34960 18386 35012
rect 21358 35000 21364 35012
rect 21319 34972 21364 35000
rect 21358 34960 21364 34972
rect 21416 34960 21422 35012
rect 23658 34932 23664 34944
rect 16908 34904 17356 34932
rect 23619 34904 23664 34932
rect 16908 34892 16914 34904
rect 23658 34892 23664 34904
rect 23716 34892 23722 34944
rect 23860 34932 23888 35031
rect 26234 35028 26240 35080
rect 26292 35028 26298 35080
rect 25130 35000 25136 35012
rect 25091 34972 25136 35000
rect 25130 34960 25136 34972
rect 25188 34960 25194 35012
rect 25222 34932 25228 34944
rect 23860 34904 25228 34932
rect 25222 34892 25228 34904
rect 25280 34892 25286 34944
rect 26602 34932 26608 34944
rect 26563 34904 26608 34932
rect 26602 34892 26608 34904
rect 26660 34892 26666 34944
rect 26712 34932 26740 35244
rect 27338 35232 27344 35244
rect 27396 35232 27402 35284
rect 28534 35232 28540 35284
rect 28592 35272 28598 35284
rect 29549 35275 29607 35281
rect 29549 35272 29561 35275
rect 28592 35244 29561 35272
rect 28592 35232 28598 35244
rect 29549 35241 29561 35244
rect 29595 35241 29607 35275
rect 32398 35272 32404 35284
rect 32359 35244 32404 35272
rect 29549 35235 29607 35241
rect 32398 35232 32404 35244
rect 32456 35232 32462 35284
rect 36722 35232 36728 35284
rect 36780 35272 36786 35284
rect 37918 35272 37924 35284
rect 36780 35244 37924 35272
rect 36780 35232 36786 35244
rect 37918 35232 37924 35244
rect 37976 35232 37982 35284
rect 28813 35207 28871 35213
rect 28813 35173 28825 35207
rect 28859 35173 28871 35207
rect 28813 35167 28871 35173
rect 27709 35139 27767 35145
rect 27709 35105 27721 35139
rect 27755 35136 27767 35139
rect 28828 35136 28856 35167
rect 31021 35139 31079 35145
rect 31021 35136 31033 35139
rect 27755 35108 28672 35136
rect 28828 35108 31033 35136
rect 27755 35105 27767 35108
rect 27709 35099 27767 35105
rect 27522 35068 27528 35080
rect 27483 35040 27528 35068
rect 27522 35028 27528 35040
rect 27580 35028 27586 35080
rect 28258 35068 28264 35080
rect 28219 35040 28264 35068
rect 28258 35028 28264 35040
rect 28316 35028 28322 35080
rect 28534 35068 28540 35080
rect 28495 35040 28540 35068
rect 28534 35028 28540 35040
rect 28592 35028 28598 35080
rect 28644 35077 28672 35108
rect 31021 35105 31033 35108
rect 31067 35105 31079 35139
rect 37182 35136 37188 35148
rect 37143 35108 37188 35136
rect 31021 35099 31079 35105
rect 37182 35096 37188 35108
rect 37240 35096 37246 35148
rect 28629 35071 28687 35077
rect 28629 35037 28641 35071
rect 28675 35068 28687 35071
rect 28994 35068 29000 35080
rect 28675 35040 29000 35068
rect 28675 35037 28687 35040
rect 28629 35031 28687 35037
rect 28994 35028 29000 35040
rect 29052 35028 29058 35080
rect 29914 35028 29920 35080
rect 29972 35028 29978 35080
rect 31294 35028 31300 35080
rect 31352 35068 31358 35080
rect 35805 35071 35863 35077
rect 31352 35040 31397 35068
rect 31352 35028 31358 35040
rect 35805 35037 35817 35071
rect 35851 35068 35863 35071
rect 36722 35068 36728 35080
rect 35851 35040 36728 35068
rect 35851 35037 35863 35040
rect 35805 35031 35863 35037
rect 36722 35028 36728 35040
rect 36780 35028 36786 35080
rect 38102 35028 38108 35080
rect 38160 35068 38166 35080
rect 38160 35040 38205 35068
rect 38160 35028 38166 35040
rect 28442 35000 28448 35012
rect 28403 34972 28448 35000
rect 28442 34960 28448 34972
rect 28500 34960 28506 35012
rect 37550 34960 37556 35012
rect 37608 35000 37614 35012
rect 37921 35003 37979 35009
rect 37921 35000 37933 35003
rect 37608 34972 37933 35000
rect 37608 34960 37614 34972
rect 37921 34969 37933 34972
rect 37967 34969 37979 35003
rect 37921 34963 37979 34969
rect 31386 34932 31392 34944
rect 26712 34904 31392 34932
rect 31386 34892 31392 34904
rect 31444 34892 31450 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2222 34728 2228 34740
rect 2183 34700 2228 34728
rect 2222 34688 2228 34700
rect 2280 34688 2286 34740
rect 2866 34728 2872 34740
rect 2827 34700 2872 34728
rect 2866 34688 2872 34700
rect 2924 34688 2930 34740
rect 10778 34728 10784 34740
rect 10739 34700 10784 34728
rect 10778 34688 10784 34700
rect 10836 34688 10842 34740
rect 12710 34728 12716 34740
rect 12406 34700 12716 34728
rect 4706 34660 4712 34672
rect 2976 34632 4712 34660
rect 1673 34595 1731 34601
rect 1673 34561 1685 34595
rect 1719 34592 1731 34595
rect 1762 34592 1768 34604
rect 1719 34564 1768 34592
rect 1719 34561 1731 34564
rect 1673 34555 1731 34561
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 2314 34592 2320 34604
rect 2275 34564 2320 34592
rect 2314 34552 2320 34564
rect 2372 34552 2378 34604
rect 2976 34601 3004 34632
rect 4706 34620 4712 34632
rect 4764 34620 4770 34672
rect 10594 34620 10600 34672
rect 10652 34660 10658 34672
rect 11517 34663 11575 34669
rect 11517 34660 11529 34663
rect 10652 34632 11529 34660
rect 10652 34620 10658 34632
rect 11517 34629 11529 34632
rect 11563 34629 11575 34663
rect 11882 34660 11888 34672
rect 11843 34632 11888 34660
rect 11517 34623 11575 34629
rect 11882 34620 11888 34632
rect 11940 34620 11946 34672
rect 12023 34663 12081 34669
rect 12023 34629 12035 34663
rect 12069 34660 12081 34663
rect 12406 34660 12434 34700
rect 12710 34688 12716 34700
rect 12768 34688 12774 34740
rect 12989 34731 13047 34737
rect 12989 34697 13001 34731
rect 13035 34728 13047 34731
rect 14182 34728 14188 34740
rect 13035 34700 14188 34728
rect 13035 34697 13047 34700
rect 12989 34691 13047 34697
rect 14182 34688 14188 34700
rect 14240 34688 14246 34740
rect 15102 34728 15108 34740
rect 15063 34700 15108 34728
rect 15102 34688 15108 34700
rect 15160 34688 15166 34740
rect 15304 34700 15608 34728
rect 12069 34632 12434 34660
rect 12621 34663 12679 34669
rect 12069 34629 12081 34632
rect 12023 34623 12081 34629
rect 12621 34629 12633 34663
rect 12667 34629 12679 34663
rect 12621 34623 12679 34629
rect 12837 34663 12895 34669
rect 12837 34629 12849 34663
rect 12883 34660 12895 34663
rect 13906 34660 13912 34672
rect 12883 34632 13912 34660
rect 12883 34629 12895 34632
rect 12837 34623 12895 34629
rect 2961 34595 3019 34601
rect 2961 34561 2973 34595
rect 3007 34561 3019 34595
rect 2961 34555 3019 34561
rect 9858 34552 9864 34604
rect 9916 34552 9922 34604
rect 10873 34595 10931 34601
rect 10873 34561 10885 34595
rect 10919 34592 10931 34595
rect 11698 34592 11704 34604
rect 10919 34564 11008 34592
rect 11659 34564 11704 34592
rect 10919 34561 10931 34564
rect 10873 34555 10931 34561
rect 3602 34524 3608 34536
rect 3563 34496 3608 34524
rect 3602 34484 3608 34496
rect 3660 34484 3666 34536
rect 3786 34524 3792 34536
rect 3747 34496 3792 34524
rect 3786 34484 3792 34496
rect 3844 34484 3850 34536
rect 3970 34484 3976 34536
rect 4028 34524 4034 34536
rect 4157 34527 4215 34533
rect 4157 34524 4169 34527
rect 4028 34496 4169 34524
rect 4028 34484 4034 34496
rect 4157 34493 4169 34496
rect 4203 34493 4215 34527
rect 8478 34524 8484 34536
rect 8439 34496 8484 34524
rect 4157 34487 4215 34493
rect 8478 34484 8484 34496
rect 8536 34484 8542 34536
rect 9950 34416 9956 34468
rect 10008 34456 10014 34468
rect 10980 34456 11008 34564
rect 11698 34552 11704 34564
rect 11756 34552 11762 34604
rect 11793 34595 11851 34601
rect 11793 34561 11805 34595
rect 11839 34561 11851 34595
rect 11793 34555 11851 34561
rect 11054 34484 11060 34536
rect 11112 34524 11118 34536
rect 11808 34524 11836 34555
rect 12158 34552 12164 34604
rect 12216 34592 12222 34604
rect 12636 34592 12664 34623
rect 13906 34620 13912 34632
rect 13964 34620 13970 34672
rect 14090 34620 14096 34672
rect 14148 34660 14154 34672
rect 14461 34663 14519 34669
rect 14461 34660 14473 34663
rect 14148 34632 14473 34660
rect 14148 34620 14154 34632
rect 14461 34629 14473 34632
rect 14507 34660 14519 34663
rect 15304 34660 15332 34700
rect 14507 34632 15332 34660
rect 14507 34629 14519 34632
rect 14461 34623 14519 34629
rect 12216 34564 12664 34592
rect 13924 34592 13952 34620
rect 14001 34595 14059 34601
rect 14001 34592 14013 34595
rect 13924 34564 14013 34592
rect 12216 34552 12222 34564
rect 14001 34561 14013 34564
rect 14047 34592 14059 34595
rect 14274 34592 14280 34604
rect 14047 34564 14280 34592
rect 14047 34561 14059 34564
rect 14001 34555 14059 34561
rect 14274 34552 14280 34564
rect 14332 34552 14338 34604
rect 15378 34552 15384 34604
rect 15436 34592 15442 34604
rect 15580 34601 15608 34700
rect 16206 34688 16212 34740
rect 16264 34728 16270 34740
rect 17129 34731 17187 34737
rect 17129 34728 17141 34731
rect 16264 34700 17141 34728
rect 16264 34688 16270 34700
rect 17129 34697 17141 34700
rect 17175 34697 17187 34731
rect 17129 34691 17187 34697
rect 17144 34660 17172 34691
rect 17402 34688 17408 34740
rect 17460 34688 17466 34740
rect 17957 34731 18015 34737
rect 17957 34697 17969 34731
rect 18003 34697 18015 34731
rect 17957 34691 18015 34697
rect 17420 34660 17448 34688
rect 17144 34632 17816 34660
rect 15565 34595 15623 34601
rect 15436 34564 15481 34592
rect 15436 34552 15442 34564
rect 15565 34561 15577 34595
rect 15611 34561 15623 34595
rect 15565 34555 15623 34561
rect 17221 34595 17279 34601
rect 17221 34561 17233 34595
rect 17267 34592 17279 34595
rect 17402 34592 17408 34604
rect 17267 34564 17408 34592
rect 17267 34561 17279 34564
rect 17221 34555 17279 34561
rect 17402 34552 17408 34564
rect 17460 34552 17466 34604
rect 17788 34601 17816 34632
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34561 17831 34595
rect 17773 34555 17831 34561
rect 11112 34496 11836 34524
rect 11112 34484 11118 34496
rect 12066 34484 12072 34536
rect 12124 34484 12130 34536
rect 14185 34527 14243 34533
rect 14185 34493 14197 34527
rect 14231 34524 14243 34527
rect 15286 34524 15292 34536
rect 14231 34496 15148 34524
rect 15247 34496 15292 34524
rect 14231 34493 14243 34496
rect 14185 34487 14243 34493
rect 12084 34456 12112 34484
rect 13170 34456 13176 34468
rect 10008 34428 13176 34456
rect 10008 34416 10014 34428
rect 13170 34416 13176 34428
rect 13228 34416 13234 34468
rect 13538 34416 13544 34468
rect 13596 34456 13602 34468
rect 15120 34456 15148 34496
rect 15286 34484 15292 34496
rect 15344 34484 15350 34536
rect 15470 34484 15476 34536
rect 15528 34524 15534 34536
rect 17972 34524 18000 34691
rect 21910 34688 21916 34740
rect 21968 34728 21974 34740
rect 22281 34731 22339 34737
rect 22281 34728 22293 34731
rect 21968 34700 22293 34728
rect 21968 34688 21974 34700
rect 22281 34697 22293 34700
rect 22327 34697 22339 34731
rect 24854 34728 24860 34740
rect 22281 34691 22339 34697
rect 23400 34700 24860 34728
rect 20714 34620 20720 34672
rect 20772 34660 20778 34672
rect 23400 34660 23428 34700
rect 24854 34688 24860 34700
rect 24912 34688 24918 34740
rect 25498 34728 25504 34740
rect 25459 34700 25504 34728
rect 25498 34688 25504 34700
rect 25556 34688 25562 34740
rect 27985 34731 28043 34737
rect 27985 34697 27997 34731
rect 28031 34728 28043 34731
rect 28626 34728 28632 34740
rect 28031 34700 28632 34728
rect 28031 34697 28043 34700
rect 27985 34691 28043 34697
rect 28626 34688 28632 34700
rect 28684 34688 28690 34740
rect 28994 34728 29000 34740
rect 28955 34700 29000 34728
rect 28994 34688 29000 34700
rect 29052 34688 29058 34740
rect 31110 34728 31116 34740
rect 29932 34700 31116 34728
rect 20772 34632 21220 34660
rect 20772 34620 20778 34632
rect 18966 34592 18972 34604
rect 18927 34564 18972 34592
rect 18966 34552 18972 34564
rect 19024 34552 19030 34604
rect 20073 34595 20131 34601
rect 20073 34561 20085 34595
rect 20119 34592 20131 34595
rect 20806 34592 20812 34604
rect 20119 34564 20812 34592
rect 20119 34561 20131 34564
rect 20073 34555 20131 34561
rect 20806 34552 20812 34564
rect 20864 34552 20870 34604
rect 21192 34601 21220 34632
rect 23308 34632 23428 34660
rect 23569 34663 23627 34669
rect 21177 34595 21235 34601
rect 21177 34561 21189 34595
rect 21223 34561 21235 34595
rect 22462 34592 22468 34604
rect 22423 34564 22468 34592
rect 21177 34555 21235 34561
rect 22462 34552 22468 34564
rect 22520 34552 22526 34604
rect 23308 34601 23336 34632
rect 23569 34629 23581 34663
rect 23615 34660 23627 34663
rect 23658 34660 23664 34672
rect 23615 34632 23664 34660
rect 23615 34629 23627 34632
rect 23569 34623 23627 34629
rect 23658 34620 23664 34632
rect 23716 34620 23722 34672
rect 25038 34660 25044 34672
rect 24794 34632 25044 34660
rect 25038 34620 25044 34632
rect 25096 34620 25102 34672
rect 26878 34660 26884 34672
rect 25148 34632 26884 34660
rect 23293 34595 23351 34601
rect 23293 34561 23305 34595
rect 23339 34561 23351 34595
rect 25148 34592 25176 34632
rect 26878 34620 26884 34632
rect 26936 34620 26942 34672
rect 27157 34663 27215 34669
rect 27157 34629 27169 34663
rect 27203 34629 27215 34663
rect 27157 34623 27215 34629
rect 27373 34663 27431 34669
rect 27373 34629 27385 34663
rect 27419 34660 27431 34663
rect 27706 34660 27712 34672
rect 27419 34632 27712 34660
rect 27419 34629 27431 34632
rect 27373 34623 27431 34629
rect 25866 34592 25872 34604
rect 23293 34555 23351 34561
rect 24872 34564 25176 34592
rect 25827 34564 25872 34592
rect 18874 34524 18880 34536
rect 15528 34496 15573 34524
rect 16500 34496 18880 34524
rect 15528 34484 15534 34496
rect 15194 34456 15200 34468
rect 13596 34428 14412 34456
rect 15120 34428 15200 34456
rect 13596 34416 13602 34428
rect 14384 34400 14412 34428
rect 15194 34416 15200 34428
rect 15252 34416 15258 34468
rect 15562 34416 15568 34468
rect 15620 34456 15626 34468
rect 16500 34456 16528 34496
rect 18874 34484 18880 34496
rect 18932 34484 18938 34536
rect 20898 34524 20904 34536
rect 20859 34496 20904 34524
rect 20898 34484 20904 34496
rect 20956 34524 20962 34536
rect 21542 34524 21548 34536
rect 20956 34496 21548 34524
rect 20956 34484 20962 34496
rect 21542 34484 21548 34496
rect 21600 34524 21606 34536
rect 24872 34524 24900 34564
rect 25866 34552 25872 34564
rect 25924 34552 25930 34604
rect 27172 34592 27200 34623
rect 27706 34620 27712 34632
rect 27764 34620 27770 34672
rect 28534 34660 28540 34672
rect 27816 34632 28396 34660
rect 28495 34632 28540 34660
rect 27816 34592 27844 34632
rect 28166 34592 28172 34604
rect 27172 34564 27844 34592
rect 28127 34564 28172 34592
rect 28166 34552 28172 34564
rect 28224 34552 28230 34604
rect 28368 34601 28396 34632
rect 28534 34620 28540 34632
rect 28592 34620 28598 34672
rect 29932 34660 29960 34700
rect 31110 34688 31116 34700
rect 31168 34688 31174 34740
rect 31386 34688 31392 34740
rect 31444 34728 31450 34740
rect 37550 34728 37556 34740
rect 31444 34700 36860 34728
rect 37511 34700 37556 34728
rect 31444 34688 31450 34700
rect 32217 34663 32275 34669
rect 32217 34660 32229 34663
rect 29840 34632 29960 34660
rect 31326 34632 32229 34660
rect 28261 34595 28319 34601
rect 28261 34561 28273 34595
rect 28307 34561 28319 34595
rect 28261 34555 28319 34561
rect 28353 34595 28411 34601
rect 28353 34561 28365 34595
rect 28399 34592 28411 34595
rect 28718 34592 28724 34604
rect 28399 34564 28724 34592
rect 28399 34561 28411 34564
rect 28353 34555 28411 34561
rect 25038 34524 25044 34536
rect 21600 34496 24900 34524
rect 24999 34496 25044 34524
rect 21600 34484 21606 34496
rect 25038 34484 25044 34496
rect 25096 34484 25102 34536
rect 25958 34524 25964 34536
rect 25919 34496 25964 34524
rect 25958 34484 25964 34496
rect 26016 34484 26022 34536
rect 26145 34527 26203 34533
rect 26145 34493 26157 34527
rect 26191 34524 26203 34527
rect 26602 34524 26608 34536
rect 26191 34496 26608 34524
rect 26191 34493 26203 34496
rect 26145 34487 26203 34493
rect 26602 34484 26608 34496
rect 26660 34484 26666 34536
rect 28276 34524 28304 34555
rect 28718 34552 28724 34564
rect 28776 34552 28782 34604
rect 28810 34552 28816 34604
rect 28868 34592 28874 34604
rect 29840 34601 29868 34632
rect 32217 34629 32229 34632
rect 32263 34629 32275 34663
rect 36538 34660 36544 34672
rect 36499 34632 36544 34660
rect 32217 34623 32275 34629
rect 36538 34620 36544 34632
rect 36596 34620 36602 34672
rect 36832 34660 36860 34700
rect 37550 34688 37556 34700
rect 37608 34688 37614 34740
rect 36832 34632 37504 34660
rect 29273 34595 29331 34601
rect 29273 34592 29285 34595
rect 28868 34564 29285 34592
rect 28868 34552 28874 34564
rect 29273 34561 29285 34564
rect 29319 34561 29331 34595
rect 29273 34555 29331 34561
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 32309 34595 32367 34601
rect 32309 34561 32321 34595
rect 32355 34592 32367 34595
rect 32398 34592 32404 34604
rect 32355 34564 32404 34592
rect 32355 34561 32367 34564
rect 32309 34555 32367 34561
rect 32398 34552 32404 34564
rect 32456 34552 32462 34604
rect 33410 34592 33416 34604
rect 33371 34564 33416 34592
rect 33410 34552 33416 34564
rect 33468 34592 33474 34604
rect 34698 34592 34704 34604
rect 33468 34564 34704 34592
rect 33468 34552 33474 34564
rect 34698 34552 34704 34564
rect 34756 34552 34762 34604
rect 36722 34552 36728 34604
rect 36780 34592 36786 34604
rect 37476 34601 37504 34632
rect 37461 34595 37519 34601
rect 36780 34564 36825 34592
rect 36780 34552 36786 34564
rect 37461 34561 37473 34595
rect 37507 34592 37519 34595
rect 38286 34592 38292 34604
rect 37507 34564 38292 34592
rect 37507 34561 37519 34564
rect 37461 34555 37519 34561
rect 38286 34552 38292 34564
rect 38344 34552 38350 34604
rect 27356 34496 28304 34524
rect 15620 34428 16528 34456
rect 15620 34416 15626 34428
rect 16758 34416 16764 34468
rect 16816 34456 16822 34468
rect 16816 34428 22094 34456
rect 16816 34416 16822 34428
rect 8744 34391 8802 34397
rect 8744 34357 8756 34391
rect 8790 34388 8802 34391
rect 10134 34388 10140 34400
rect 8790 34360 10140 34388
rect 8790 34357 8802 34360
rect 8744 34351 8802 34357
rect 10134 34348 10140 34360
rect 10192 34348 10198 34400
rect 10229 34391 10287 34397
rect 10229 34357 10241 34391
rect 10275 34388 10287 34391
rect 11974 34388 11980 34400
rect 10275 34360 11980 34388
rect 10275 34357 10287 34360
rect 10229 34351 10287 34357
rect 11974 34348 11980 34360
rect 12032 34388 12038 34400
rect 12805 34391 12863 34397
rect 12805 34388 12817 34391
rect 12032 34360 12817 34388
rect 12032 34348 12038 34360
rect 12805 34357 12817 34360
rect 12851 34357 12863 34391
rect 12805 34351 12863 34357
rect 13817 34391 13875 34397
rect 13817 34357 13829 34391
rect 13863 34388 13875 34391
rect 13906 34388 13912 34400
rect 13863 34360 13912 34388
rect 13863 34357 13875 34360
rect 13817 34351 13875 34357
rect 13906 34348 13912 34360
rect 13964 34348 13970 34400
rect 14366 34388 14372 34400
rect 14327 34360 14372 34388
rect 14366 34348 14372 34360
rect 14424 34348 14430 34400
rect 15102 34348 15108 34400
rect 15160 34388 15166 34400
rect 17862 34388 17868 34400
rect 15160 34360 17868 34388
rect 15160 34348 15166 34360
rect 17862 34348 17868 34360
rect 17920 34348 17926 34400
rect 18506 34348 18512 34400
rect 18564 34388 18570 34400
rect 18877 34391 18935 34397
rect 18877 34388 18889 34391
rect 18564 34360 18889 34388
rect 18564 34348 18570 34360
rect 18877 34357 18889 34360
rect 18923 34357 18935 34391
rect 19978 34388 19984 34400
rect 19939 34360 19984 34388
rect 18877 34351 18935 34357
rect 19978 34348 19984 34360
rect 20036 34348 20042 34400
rect 22066 34388 22094 34428
rect 25774 34388 25780 34400
rect 22066 34360 25780 34388
rect 25774 34348 25780 34360
rect 25832 34348 25838 34400
rect 26620 34388 26648 34484
rect 27356 34400 27384 34496
rect 28534 34484 28540 34536
rect 28592 34524 28598 34536
rect 28828 34524 28856 34552
rect 28994 34524 29000 34536
rect 28592 34496 28856 34524
rect 28955 34496 29000 34524
rect 28592 34484 28598 34496
rect 28994 34484 29000 34496
rect 29052 34484 29058 34536
rect 33778 34524 33784 34536
rect 33739 34496 33784 34524
rect 33778 34484 33784 34496
rect 33836 34484 33842 34536
rect 35802 34524 35808 34536
rect 35763 34496 35808 34524
rect 35802 34484 35808 34496
rect 35860 34484 35866 34536
rect 27525 34459 27583 34465
rect 27525 34425 27537 34459
rect 27571 34456 27583 34459
rect 28258 34456 28264 34468
rect 27571 34428 28264 34456
rect 27571 34425 27583 34428
rect 27525 34419 27583 34425
rect 28258 34416 28264 34428
rect 28316 34456 28322 34468
rect 29181 34459 29239 34465
rect 29181 34456 29193 34459
rect 28316 34428 29193 34456
rect 28316 34416 28322 34428
rect 29181 34425 29193 34428
rect 29227 34425 29239 34459
rect 29181 34419 29239 34425
rect 27338 34388 27344 34400
rect 26620 34360 27344 34388
rect 27338 34348 27344 34360
rect 27396 34348 27402 34400
rect 30088 34391 30146 34397
rect 30088 34357 30100 34391
rect 30134 34388 30146 34391
rect 30650 34388 30656 34400
rect 30134 34360 30656 34388
rect 30134 34357 30146 34360
rect 30088 34351 30146 34357
rect 30650 34348 30656 34360
rect 30708 34348 30714 34400
rect 30742 34348 30748 34400
rect 30800 34388 30806 34400
rect 31573 34391 31631 34397
rect 31573 34388 31585 34391
rect 30800 34360 31585 34388
rect 30800 34348 30806 34360
rect 31573 34357 31585 34360
rect 31619 34357 31631 34391
rect 31573 34351 31631 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1949 34187 2007 34193
rect 1949 34153 1961 34187
rect 1995 34184 2007 34187
rect 3234 34184 3240 34196
rect 1995 34156 3240 34184
rect 1995 34153 2007 34156
rect 1949 34147 2007 34153
rect 3234 34144 3240 34156
rect 3292 34144 3298 34196
rect 3786 34144 3792 34196
rect 3844 34184 3850 34196
rect 3881 34187 3939 34193
rect 3881 34184 3893 34187
rect 3844 34156 3893 34184
rect 3844 34144 3850 34156
rect 3881 34153 3893 34156
rect 3927 34153 3939 34187
rect 5626 34184 5632 34196
rect 3881 34147 3939 34153
rect 4356 34156 5632 34184
rect 2593 34119 2651 34125
rect 2593 34085 2605 34119
rect 2639 34116 2651 34119
rect 3418 34116 3424 34128
rect 2639 34088 3424 34116
rect 2639 34085 2651 34088
rect 2593 34079 2651 34085
rect 3418 34076 3424 34088
rect 3476 34076 3482 34128
rect 3237 34051 3295 34057
rect 3237 34017 3249 34051
rect 3283 34048 3295 34051
rect 4356 34048 4384 34156
rect 5626 34144 5632 34156
rect 5684 34144 5690 34196
rect 5994 34144 6000 34196
rect 6052 34184 6058 34196
rect 9858 34184 9864 34196
rect 6052 34156 6914 34184
rect 9819 34156 9864 34184
rect 6052 34144 6058 34156
rect 5718 34116 5724 34128
rect 3283 34020 4384 34048
rect 4448 34088 5724 34116
rect 3283 34017 3295 34020
rect 3237 34011 3295 34017
rect 4448 33989 4476 34088
rect 5718 34076 5724 34088
rect 5776 34076 5782 34128
rect 6886 34116 6914 34156
rect 9858 34144 9864 34156
rect 9916 34144 9922 34196
rect 10134 34144 10140 34196
rect 10192 34184 10198 34196
rect 11701 34187 11759 34193
rect 11701 34184 11713 34187
rect 10192 34156 11713 34184
rect 10192 34144 10198 34156
rect 11701 34153 11713 34156
rect 11747 34153 11759 34187
rect 11701 34147 11759 34153
rect 11790 34144 11796 34196
rect 11848 34184 11854 34196
rect 14277 34187 14335 34193
rect 11848 34156 14228 34184
rect 11848 34144 11854 34156
rect 14200 34116 14228 34156
rect 14277 34153 14289 34187
rect 14323 34184 14335 34187
rect 14458 34184 14464 34196
rect 14323 34156 14464 34184
rect 14323 34153 14335 34156
rect 14277 34147 14335 34153
rect 14458 34144 14464 34156
rect 14516 34144 14522 34196
rect 16206 34184 16212 34196
rect 14568 34156 16212 34184
rect 14568 34116 14596 34156
rect 16206 34144 16212 34156
rect 16264 34144 16270 34196
rect 16298 34144 16304 34196
rect 16356 34184 16362 34196
rect 17129 34187 17187 34193
rect 17129 34184 17141 34187
rect 16356 34156 17141 34184
rect 16356 34144 16362 34156
rect 17129 34153 17141 34156
rect 17175 34153 17187 34187
rect 17129 34147 17187 34153
rect 17862 34144 17868 34196
rect 17920 34184 17926 34196
rect 20990 34184 20996 34196
rect 17920 34156 20996 34184
rect 17920 34144 17926 34156
rect 20990 34144 20996 34156
rect 21048 34144 21054 34196
rect 25222 34184 25228 34196
rect 25183 34156 25228 34184
rect 25222 34144 25228 34156
rect 25280 34144 25286 34196
rect 28994 34184 29000 34196
rect 25332 34156 29000 34184
rect 6886 34088 14136 34116
rect 14200 34088 14596 34116
rect 10965 34051 11023 34057
rect 10965 34017 10977 34051
rect 11011 34048 11023 34051
rect 11146 34048 11152 34060
rect 11011 34020 11152 34048
rect 11011 34017 11023 34020
rect 10965 34011 11023 34017
rect 11146 34008 11152 34020
rect 11204 34008 11210 34060
rect 11241 34051 11299 34057
rect 11241 34017 11253 34051
rect 11287 34048 11299 34051
rect 13814 34048 13820 34060
rect 11287 34020 12296 34048
rect 11287 34017 11299 34020
rect 11241 34011 11299 34017
rect 3973 33983 4031 33989
rect 3973 33949 3985 33983
rect 4019 33949 4031 33983
rect 3973 33943 4031 33949
rect 4433 33983 4491 33989
rect 4433 33949 4445 33983
rect 4479 33949 4491 33983
rect 4433 33943 4491 33949
rect 5353 33983 5411 33989
rect 5353 33949 5365 33983
rect 5399 33980 5411 33983
rect 5810 33980 5816 33992
rect 5399 33952 5816 33980
rect 5399 33949 5411 33952
rect 5353 33943 5411 33949
rect 3988 33912 4016 33943
rect 5258 33912 5264 33924
rect 3988 33884 5264 33912
rect 5258 33872 5264 33884
rect 5316 33872 5322 33924
rect 4617 33847 4675 33853
rect 4617 33813 4629 33847
rect 4663 33844 4675 33847
rect 5368 33844 5396 33943
rect 5810 33940 5816 33952
rect 5868 33980 5874 33992
rect 6641 33983 6699 33989
rect 6641 33980 6653 33983
rect 5868 33952 6653 33980
rect 5868 33940 5874 33952
rect 6641 33949 6653 33952
rect 6687 33949 6699 33983
rect 9950 33980 9956 33992
rect 9911 33952 9956 33980
rect 6641 33943 6699 33949
rect 9950 33940 9956 33952
rect 10008 33940 10014 33992
rect 10873 33983 10931 33989
rect 10873 33949 10885 33983
rect 10919 33949 10931 33983
rect 10873 33943 10931 33949
rect 5994 33912 6000 33924
rect 5955 33884 6000 33912
rect 5994 33872 6000 33884
rect 6052 33872 6058 33924
rect 7466 33912 7472 33924
rect 7427 33884 7472 33912
rect 7466 33872 7472 33884
rect 7524 33872 7530 33924
rect 10888 33912 10916 33943
rect 11790 33940 11796 33992
rect 11848 33980 11854 33992
rect 11885 33983 11943 33989
rect 11885 33980 11897 33983
rect 11848 33952 11897 33980
rect 11848 33940 11854 33952
rect 11885 33949 11897 33952
rect 11931 33949 11943 33983
rect 11885 33943 11943 33949
rect 11974 33940 11980 33992
rect 12032 33980 12038 33992
rect 12268 33989 12296 34020
rect 13096 34020 13820 34048
rect 12253 33983 12311 33989
rect 12032 33952 12077 33980
rect 12032 33940 12038 33952
rect 12253 33949 12265 33983
rect 12299 33949 12311 33983
rect 12253 33943 12311 33949
rect 12526 33940 12532 33992
rect 12584 33980 12590 33992
rect 13096 33989 13124 34020
rect 13814 34008 13820 34020
rect 13872 34008 13878 34060
rect 14108 34048 14136 34088
rect 17034 34076 17040 34128
rect 17092 34116 17098 34128
rect 18417 34119 18475 34125
rect 18417 34116 18429 34119
rect 17092 34088 18429 34116
rect 17092 34076 17098 34088
rect 18417 34085 18429 34088
rect 18463 34085 18475 34119
rect 18417 34079 18475 34085
rect 24118 34076 24124 34128
rect 24176 34116 24182 34128
rect 25332 34116 25360 34156
rect 28994 34144 29000 34156
rect 29052 34144 29058 34196
rect 29914 34184 29920 34196
rect 29875 34156 29920 34184
rect 29914 34144 29920 34156
rect 29972 34144 29978 34196
rect 24176 34088 25360 34116
rect 24176 34076 24182 34088
rect 26970 34076 26976 34128
rect 27028 34116 27034 34128
rect 30098 34116 30104 34128
rect 27028 34088 30104 34116
rect 27028 34076 27034 34088
rect 15102 34048 15108 34060
rect 14108 34020 15108 34048
rect 15102 34008 15108 34020
rect 15160 34008 15166 34060
rect 15378 34048 15384 34060
rect 15291 34020 15384 34048
rect 15378 34008 15384 34020
rect 15436 34048 15442 34060
rect 16390 34048 16396 34060
rect 15436 34020 16396 34048
rect 15436 34008 15442 34020
rect 16390 34008 16396 34020
rect 16448 34008 16454 34060
rect 18325 34051 18383 34057
rect 18325 34017 18337 34051
rect 18371 34048 18383 34051
rect 18598 34048 18604 34060
rect 18371 34020 18604 34048
rect 18371 34017 18383 34020
rect 18325 34011 18383 34017
rect 18598 34008 18604 34020
rect 18656 34008 18662 34060
rect 18693 34051 18751 34057
rect 18693 34017 18705 34051
rect 18739 34048 18751 34051
rect 20717 34051 20775 34057
rect 20717 34048 20729 34051
rect 18739 34020 20729 34048
rect 18739 34017 18751 34020
rect 18693 34011 18751 34017
rect 20717 34017 20729 34020
rect 20763 34017 20775 34051
rect 21910 34048 21916 34060
rect 21871 34020 21916 34048
rect 20717 34011 20775 34017
rect 21910 34008 21916 34020
rect 21968 34008 21974 34060
rect 23382 34008 23388 34060
rect 23440 34048 23446 34060
rect 25593 34051 25651 34057
rect 25593 34048 25605 34051
rect 23440 34020 25605 34048
rect 23440 34008 23446 34020
rect 25593 34017 25605 34020
rect 25639 34017 25651 34051
rect 25593 34011 25651 34017
rect 27338 34008 27344 34060
rect 27396 34048 27402 34060
rect 27893 34051 27951 34057
rect 27893 34048 27905 34051
rect 27396 34020 27905 34048
rect 27396 34008 27402 34020
rect 27893 34017 27905 34020
rect 27939 34017 27951 34051
rect 27893 34011 27951 34017
rect 27985 34051 28043 34057
rect 27985 34017 27997 34051
rect 28031 34048 28043 34051
rect 28718 34048 28724 34060
rect 28031 34020 28724 34048
rect 28031 34017 28043 34020
rect 27985 34011 28043 34017
rect 28718 34008 28724 34020
rect 28776 34008 28782 34060
rect 12989 33983 13047 33989
rect 12989 33980 13001 33983
rect 12584 33952 13001 33980
rect 12584 33940 12590 33952
rect 12989 33949 13001 33952
rect 13035 33949 13047 33983
rect 12989 33943 13047 33949
rect 13081 33983 13139 33989
rect 13081 33949 13093 33983
rect 13127 33949 13139 33983
rect 13262 33980 13268 33992
rect 13223 33952 13268 33980
rect 13081 33943 13139 33949
rect 13262 33940 13268 33952
rect 13320 33940 13326 33992
rect 13357 33983 13415 33989
rect 13357 33949 13369 33983
rect 13403 33949 13415 33983
rect 18230 33980 18236 33992
rect 18191 33952 18236 33980
rect 13357 33943 13415 33949
rect 11146 33912 11152 33924
rect 10888 33884 11152 33912
rect 11146 33872 11152 33884
rect 11204 33912 11210 33924
rect 11992 33912 12020 33940
rect 11204 33884 12020 33912
rect 12069 33915 12127 33921
rect 11204 33872 11210 33884
rect 12069 33881 12081 33915
rect 12115 33912 12127 33915
rect 12618 33912 12624 33924
rect 12115 33884 12624 33912
rect 12115 33881 12127 33884
rect 12069 33875 12127 33881
rect 12618 33872 12624 33884
rect 12676 33872 12682 33924
rect 13372 33912 13400 33943
rect 18230 33940 18236 33952
rect 18288 33940 18294 33992
rect 18506 33940 18512 33992
rect 18564 33980 18570 33992
rect 18564 33952 18609 33980
rect 18564 33940 18570 33952
rect 20990 33940 20996 33992
rect 21048 33980 21054 33992
rect 21637 33983 21695 33989
rect 21637 33980 21649 33983
rect 21048 33952 21649 33980
rect 21048 33940 21054 33952
rect 21637 33949 21649 33952
rect 21683 33949 21695 33983
rect 21637 33943 21695 33949
rect 24210 33940 24216 33992
rect 24268 33980 24274 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 24268 33952 24593 33980
rect 24268 33940 24274 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 24670 33940 24676 33992
rect 24728 33980 24734 33992
rect 24728 33952 24773 33980
rect 24728 33940 24734 33952
rect 24946 33940 24952 33992
rect 25004 33980 25010 33992
rect 25409 33983 25467 33989
rect 25409 33980 25421 33983
rect 25004 33952 25421 33980
rect 25004 33940 25010 33952
rect 25409 33949 25421 33952
rect 25455 33949 25467 33983
rect 25409 33943 25467 33949
rect 25958 33940 25964 33992
rect 26016 33980 26022 33992
rect 26053 33983 26111 33989
rect 26053 33980 26065 33983
rect 26016 33952 26065 33980
rect 26016 33940 26022 33952
rect 26053 33949 26065 33952
rect 26099 33949 26111 33983
rect 26234 33980 26240 33992
rect 26195 33952 26240 33980
rect 26053 33943 26111 33949
rect 26234 33940 26240 33952
rect 26292 33940 26298 33992
rect 26421 33983 26479 33989
rect 26421 33949 26433 33983
rect 26467 33980 26479 33983
rect 27065 33983 27123 33989
rect 27065 33980 27077 33983
rect 26467 33952 27077 33980
rect 26467 33949 26479 33952
rect 26421 33943 26479 33949
rect 27065 33949 27077 33952
rect 27111 33949 27123 33983
rect 27706 33980 27712 33992
rect 27667 33952 27712 33980
rect 27065 33943 27123 33949
rect 27706 33940 27712 33952
rect 27764 33940 27770 33992
rect 29840 33989 29868 34088
rect 30098 34076 30104 34088
rect 30156 34076 30162 34128
rect 32398 34048 32404 34060
rect 30668 34020 32404 34048
rect 27801 33983 27859 33989
rect 27801 33949 27813 33983
rect 27847 33949 27859 33983
rect 27801 33943 27859 33949
rect 29825 33983 29883 33989
rect 29825 33949 29837 33983
rect 29871 33980 29883 33983
rect 29914 33980 29920 33992
rect 29871 33952 29920 33980
rect 29871 33949 29883 33952
rect 29825 33943 29883 33949
rect 12728 33884 13400 33912
rect 4663 33816 5396 33844
rect 4663 33813 4675 33816
rect 4617 33807 4675 33813
rect 10134 33804 10140 33856
rect 10192 33844 10198 33856
rect 11698 33844 11704 33856
rect 10192 33816 11704 33844
rect 10192 33804 10198 33816
rect 11698 33804 11704 33816
rect 11756 33804 11762 33856
rect 11882 33804 11888 33856
rect 11940 33844 11946 33856
rect 12728 33844 12756 33884
rect 14182 33872 14188 33924
rect 14240 33921 14246 33924
rect 14240 33915 14303 33921
rect 14240 33881 14257 33915
rect 14291 33881 14303 33915
rect 14240 33875 14303 33881
rect 14240 33872 14246 33875
rect 14366 33872 14372 33924
rect 14424 33912 14430 33924
rect 14461 33915 14519 33921
rect 14461 33912 14473 33915
rect 14424 33884 14473 33912
rect 14424 33872 14430 33884
rect 14461 33881 14473 33884
rect 14507 33881 14519 33915
rect 15654 33912 15660 33924
rect 15615 33884 15660 33912
rect 14461 33875 14519 33881
rect 15654 33872 15660 33884
rect 15712 33872 15718 33924
rect 16942 33912 16948 33924
rect 16882 33884 16948 33912
rect 16942 33872 16948 33884
rect 17000 33872 17006 33924
rect 19334 33912 19340 33924
rect 18892 33884 19340 33912
rect 11940 33816 12756 33844
rect 12805 33847 12863 33853
rect 11940 33804 11946 33816
rect 12805 33813 12817 33847
rect 12851 33844 12863 33847
rect 13078 33844 13084 33856
rect 12851 33816 13084 33844
rect 12851 33813 12863 33816
rect 12805 33807 12863 33813
rect 13078 33804 13084 33816
rect 13136 33804 13142 33856
rect 13262 33804 13268 33856
rect 13320 33844 13326 33856
rect 14093 33847 14151 33853
rect 14093 33844 14105 33847
rect 13320 33816 14105 33844
rect 13320 33804 13326 33816
rect 14093 33813 14105 33816
rect 14139 33813 14151 33847
rect 14093 33807 14151 33813
rect 15194 33804 15200 33856
rect 15252 33844 15258 33856
rect 18892 33844 18920 33884
rect 19334 33872 19340 33884
rect 19392 33872 19398 33924
rect 19978 33872 19984 33924
rect 20036 33872 20042 33924
rect 22646 33872 22652 33924
rect 22704 33872 22710 33924
rect 24688 33912 24716 33940
rect 26694 33912 26700 33924
rect 24688 33884 26700 33912
rect 26694 33872 26700 33884
rect 26752 33912 26758 33924
rect 27816 33912 27844 33943
rect 29914 33940 29920 33952
rect 29972 33940 29978 33992
rect 30558 33940 30564 33992
rect 30616 33980 30622 33992
rect 30668 33989 30696 34020
rect 32398 34008 32404 34020
rect 32456 34008 32462 34060
rect 37366 34048 37372 34060
rect 37327 34020 37372 34048
rect 37366 34008 37372 34020
rect 37424 34008 37430 34060
rect 30653 33983 30711 33989
rect 30653 33980 30665 33983
rect 30616 33952 30665 33980
rect 30616 33940 30622 33952
rect 30653 33949 30665 33952
rect 30699 33949 30711 33983
rect 30653 33943 30711 33949
rect 30926 33940 30932 33992
rect 30984 33980 30990 33992
rect 31294 33980 31300 33992
rect 30984 33952 31300 33980
rect 30984 33940 30990 33952
rect 31294 33940 31300 33952
rect 31352 33980 31358 33992
rect 32033 33983 32091 33989
rect 32033 33980 32045 33983
rect 31352 33952 32045 33980
rect 31352 33940 31358 33952
rect 32033 33949 32045 33952
rect 32079 33949 32091 33983
rect 36262 33980 36268 33992
rect 36223 33952 36268 33980
rect 32033 33943 32091 33949
rect 36262 33940 36268 33952
rect 36320 33940 36326 33992
rect 27890 33912 27896 33924
rect 26752 33884 27896 33912
rect 26752 33872 26758 33884
rect 27890 33872 27896 33884
rect 27948 33872 27954 33924
rect 32306 33912 32312 33924
rect 32267 33884 32312 33912
rect 32306 33872 32312 33884
rect 32364 33872 32370 33924
rect 33318 33872 33324 33924
rect 33376 33872 33382 33924
rect 36449 33915 36507 33921
rect 36449 33881 36461 33915
rect 36495 33912 36507 33915
rect 37366 33912 37372 33924
rect 36495 33884 37372 33912
rect 36495 33881 36507 33884
rect 36449 33875 36507 33881
rect 37366 33872 37372 33884
rect 37424 33872 37430 33924
rect 15252 33816 18920 33844
rect 15252 33804 15258 33816
rect 18966 33804 18972 33856
rect 19024 33844 19030 33856
rect 19245 33847 19303 33853
rect 19245 33844 19257 33847
rect 19024 33816 19257 33844
rect 19024 33804 19030 33816
rect 19245 33813 19257 33816
rect 19291 33813 19303 33847
rect 19245 33807 19303 33813
rect 23385 33847 23443 33853
rect 23385 33813 23397 33847
rect 23431 33844 23443 33847
rect 23474 33844 23480 33856
rect 23431 33816 23480 33844
rect 23431 33813 23443 33816
rect 23385 33807 23443 33813
rect 23474 33804 23480 33816
rect 23532 33804 23538 33856
rect 24394 33844 24400 33856
rect 24355 33816 24400 33844
rect 24394 33804 24400 33816
rect 24452 33804 24458 33856
rect 26326 33804 26332 33856
rect 26384 33844 26390 33856
rect 26881 33847 26939 33853
rect 26881 33844 26893 33847
rect 26384 33816 26893 33844
rect 26384 33804 26390 33816
rect 26881 33813 26893 33816
rect 26927 33813 26939 33847
rect 27522 33844 27528 33856
rect 27483 33816 27528 33844
rect 26881 33807 26939 33813
rect 27522 33804 27528 33816
rect 27580 33804 27586 33856
rect 30006 33804 30012 33856
rect 30064 33844 30070 33856
rect 30561 33847 30619 33853
rect 30561 33844 30573 33847
rect 30064 33816 30573 33844
rect 30064 33804 30070 33816
rect 30561 33813 30573 33816
rect 30607 33813 30619 33847
rect 30561 33807 30619 33813
rect 32122 33804 32128 33856
rect 32180 33844 32186 33856
rect 33781 33847 33839 33853
rect 33781 33844 33793 33847
rect 32180 33816 33793 33844
rect 32180 33804 32186 33816
rect 33781 33813 33793 33816
rect 33827 33813 33839 33847
rect 33781 33807 33839 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 5350 33600 5356 33652
rect 5408 33640 5414 33652
rect 14550 33640 14556 33652
rect 5408 33612 11376 33640
rect 5408 33600 5414 33612
rect 9769 33575 9827 33581
rect 9769 33541 9781 33575
rect 9815 33572 9827 33575
rect 11054 33572 11060 33584
rect 9815 33544 11060 33572
rect 9815 33541 9827 33544
rect 9769 33535 9827 33541
rect 11054 33532 11060 33544
rect 11112 33532 11118 33584
rect 2133 33507 2191 33513
rect 2133 33473 2145 33507
rect 2179 33504 2191 33507
rect 2958 33504 2964 33516
rect 2179 33476 2964 33504
rect 2179 33473 2191 33476
rect 2133 33467 2191 33473
rect 2958 33464 2964 33476
rect 3016 33464 3022 33516
rect 3602 33504 3608 33516
rect 3563 33476 3608 33504
rect 3602 33464 3608 33476
rect 3660 33464 3666 33516
rect 4985 33507 5043 33513
rect 4985 33473 4997 33507
rect 5031 33504 5043 33507
rect 5810 33504 5816 33516
rect 5031 33476 5816 33504
rect 5031 33473 5043 33476
rect 4985 33467 5043 33473
rect 5810 33464 5816 33476
rect 5868 33464 5874 33516
rect 6730 33464 6736 33516
rect 6788 33504 6794 33516
rect 8389 33507 8447 33513
rect 8389 33504 8401 33507
rect 6788 33476 8401 33504
rect 6788 33464 6794 33476
rect 8389 33473 8401 33476
rect 8435 33504 8447 33507
rect 9033 33507 9091 33513
rect 9033 33504 9045 33507
rect 8435 33476 9045 33504
rect 8435 33473 8447 33476
rect 8389 33467 8447 33473
rect 9033 33473 9045 33476
rect 9079 33473 9091 33507
rect 9033 33467 9091 33473
rect 9861 33507 9919 33513
rect 9861 33473 9873 33507
rect 9907 33504 9919 33507
rect 10226 33504 10232 33516
rect 9907 33476 10232 33504
rect 9907 33473 9919 33476
rect 9861 33467 9919 33473
rect 10226 33464 10232 33476
rect 10284 33464 10290 33516
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33504 10379 33507
rect 10597 33507 10655 33513
rect 10367 33476 10548 33504
rect 10367 33473 10379 33476
rect 10321 33467 10379 33473
rect 5350 33436 5356 33448
rect 5311 33408 5356 33436
rect 5350 33396 5356 33408
rect 5408 33396 5414 33448
rect 10413 33439 10471 33445
rect 10413 33405 10425 33439
rect 10459 33405 10471 33439
rect 10520 33436 10548 33476
rect 10597 33473 10609 33507
rect 10643 33504 10655 33507
rect 10870 33504 10876 33516
rect 10643 33476 10876 33504
rect 10643 33473 10655 33476
rect 10597 33467 10655 33473
rect 10870 33464 10876 33476
rect 10928 33464 10934 33516
rect 11146 33436 11152 33448
rect 10520 33408 11152 33436
rect 10413 33399 10471 33405
rect 3418 33328 3424 33380
rect 3476 33368 3482 33380
rect 10134 33368 10140 33380
rect 3476 33340 10140 33368
rect 3476 33328 3482 33340
rect 10134 33328 10140 33340
rect 10192 33328 10198 33380
rect 10428 33368 10456 33399
rect 11146 33396 11152 33408
rect 11204 33396 11210 33448
rect 10686 33368 10692 33380
rect 10428 33340 10692 33368
rect 10686 33328 10692 33340
rect 10744 33328 10750 33380
rect 8386 33260 8392 33312
rect 8444 33300 8450 33312
rect 8481 33303 8539 33309
rect 8481 33300 8493 33303
rect 8444 33272 8493 33300
rect 8444 33260 8450 33272
rect 8481 33269 8493 33272
rect 8527 33269 8539 33303
rect 9122 33300 9128 33312
rect 9083 33272 9128 33300
rect 8481 33263 8539 33269
rect 9122 33260 9128 33272
rect 9180 33260 9186 33312
rect 10318 33300 10324 33312
rect 10279 33272 10324 33300
rect 10318 33260 10324 33272
rect 10376 33260 10382 33312
rect 10778 33300 10784 33312
rect 10739 33272 10784 33300
rect 10778 33260 10784 33272
rect 10836 33260 10842 33312
rect 11348 33300 11376 33612
rect 11716 33612 14556 33640
rect 11716 33581 11744 33612
rect 14550 33600 14556 33612
rect 14608 33600 14614 33652
rect 15749 33643 15807 33649
rect 15749 33609 15761 33643
rect 15795 33640 15807 33643
rect 16482 33640 16488 33652
rect 15795 33612 16488 33640
rect 15795 33609 15807 33612
rect 15749 33603 15807 33609
rect 16482 33600 16488 33612
rect 16540 33600 16546 33652
rect 16945 33643 17003 33649
rect 16945 33609 16957 33643
rect 16991 33640 17003 33643
rect 17034 33640 17040 33652
rect 16991 33612 17040 33640
rect 16991 33609 17003 33612
rect 16945 33603 17003 33609
rect 17034 33600 17040 33612
rect 17092 33600 17098 33652
rect 18230 33600 18236 33652
rect 18288 33640 18294 33652
rect 18509 33643 18567 33649
rect 18509 33640 18521 33643
rect 18288 33612 18521 33640
rect 18288 33600 18294 33612
rect 18509 33609 18521 33612
rect 18555 33609 18567 33643
rect 18509 33603 18567 33609
rect 22462 33600 22468 33652
rect 22520 33640 22526 33652
rect 22925 33643 22983 33649
rect 22925 33640 22937 33643
rect 22520 33612 22937 33640
rect 22520 33600 22526 33612
rect 22925 33609 22937 33612
rect 22971 33609 22983 33643
rect 22925 33603 22983 33609
rect 23293 33643 23351 33649
rect 23293 33609 23305 33643
rect 23339 33640 23351 33643
rect 24394 33640 24400 33652
rect 23339 33612 24400 33640
rect 23339 33609 23351 33612
rect 23293 33603 23351 33609
rect 24394 33600 24400 33612
rect 24452 33600 24458 33652
rect 24946 33640 24952 33652
rect 24907 33612 24952 33640
rect 24946 33600 24952 33612
rect 25004 33600 25010 33652
rect 25777 33643 25835 33649
rect 25777 33609 25789 33643
rect 25823 33640 25835 33643
rect 25866 33640 25872 33652
rect 25823 33612 25872 33640
rect 25823 33609 25835 33612
rect 25777 33603 25835 33609
rect 25866 33600 25872 33612
rect 25924 33600 25930 33652
rect 26234 33600 26240 33652
rect 26292 33640 26298 33652
rect 27617 33643 27675 33649
rect 27617 33640 27629 33643
rect 26292 33612 27629 33640
rect 26292 33600 26298 33612
rect 27617 33609 27629 33612
rect 27663 33609 27675 33643
rect 27617 33603 27675 33609
rect 33229 33643 33287 33649
rect 33229 33609 33241 33643
rect 33275 33640 33287 33643
rect 33318 33640 33324 33652
rect 33275 33612 33324 33640
rect 33275 33609 33287 33612
rect 33229 33603 33287 33609
rect 33318 33600 33324 33612
rect 33376 33600 33382 33652
rect 37366 33640 37372 33652
rect 37327 33612 37372 33640
rect 37366 33600 37372 33612
rect 37424 33600 37430 33652
rect 11701 33575 11759 33581
rect 11701 33541 11713 33575
rect 11747 33541 11759 33575
rect 11701 33535 11759 33541
rect 11790 33532 11796 33584
rect 11848 33572 11854 33584
rect 12802 33572 12808 33584
rect 11848 33544 12808 33572
rect 11848 33532 11854 33544
rect 12802 33532 12808 33544
rect 12860 33532 12866 33584
rect 15194 33572 15200 33584
rect 14122 33544 15200 33572
rect 15194 33532 15200 33544
rect 15252 33532 15258 33584
rect 15286 33532 15292 33584
rect 15344 33532 15350 33584
rect 15381 33575 15439 33581
rect 15381 33541 15393 33575
rect 15427 33572 15439 33575
rect 17402 33572 17408 33584
rect 15427 33544 17408 33572
rect 15427 33541 15439 33544
rect 15381 33535 15439 33541
rect 17402 33532 17408 33544
rect 17460 33532 17466 33584
rect 17957 33575 18015 33581
rect 17957 33541 17969 33575
rect 18003 33572 18015 33575
rect 18414 33572 18420 33584
rect 18003 33544 18420 33572
rect 18003 33541 18015 33544
rect 17957 33535 18015 33541
rect 18414 33532 18420 33544
rect 18472 33572 18478 33584
rect 20714 33572 20720 33584
rect 18472 33544 18920 33572
rect 20562 33544 20720 33572
rect 18472 33532 18478 33544
rect 15304 33504 15332 33532
rect 18892 33513 18920 33544
rect 20714 33532 20720 33544
rect 20772 33532 20778 33584
rect 20990 33532 20996 33584
rect 21048 33572 21054 33584
rect 22189 33575 22247 33581
rect 21048 33544 21312 33572
rect 21048 33532 21054 33544
rect 21284 33513 21312 33544
rect 22189 33541 22201 33575
rect 22235 33572 22247 33575
rect 23382 33572 23388 33584
rect 22235 33544 23388 33572
rect 22235 33541 22247 33544
rect 22189 33535 22247 33541
rect 23382 33532 23388 33544
rect 23440 33532 23446 33584
rect 25222 33572 25228 33584
rect 24412 33544 25228 33572
rect 15120 33476 15332 33504
rect 17037 33507 17095 33513
rect 12342 33436 12348 33448
rect 11532 33408 12348 33436
rect 11532 33380 11560 33408
rect 12342 33396 12348 33408
rect 12400 33436 12406 33448
rect 12621 33439 12679 33445
rect 12621 33436 12633 33439
rect 12400 33408 12633 33436
rect 12400 33396 12406 33408
rect 12621 33405 12633 33408
rect 12667 33405 12679 33439
rect 12894 33436 12900 33448
rect 12855 33408 12900 33436
rect 12621 33399 12679 33405
rect 12894 33396 12900 33408
rect 12952 33396 12958 33448
rect 13354 33396 13360 33448
rect 13412 33436 13418 33448
rect 13412 33408 13952 33436
rect 13412 33396 13418 33408
rect 11514 33368 11520 33380
rect 11475 33340 11520 33368
rect 11514 33328 11520 33340
rect 11572 33328 11578 33380
rect 13924 33368 13952 33408
rect 14274 33396 14280 33448
rect 14332 33436 14338 33448
rect 15120 33445 15148 33476
rect 17037 33473 17049 33507
rect 17083 33473 17095 33507
rect 17037 33467 17095 33473
rect 18049 33507 18107 33513
rect 18049 33473 18061 33507
rect 18095 33504 18107 33507
rect 18877 33507 18935 33513
rect 18095 33476 18736 33504
rect 18095 33473 18107 33476
rect 18049 33467 18107 33473
rect 14369 33439 14427 33445
rect 14369 33436 14381 33439
rect 14332 33408 14381 33436
rect 14332 33396 14338 33408
rect 14369 33405 14381 33408
rect 14415 33405 14427 33439
rect 14369 33399 14427 33405
rect 15105 33439 15163 33445
rect 15105 33405 15117 33439
rect 15151 33405 15163 33439
rect 15286 33436 15292 33448
rect 15247 33408 15292 33436
rect 15105 33399 15163 33405
rect 15286 33396 15292 33408
rect 15344 33396 15350 33448
rect 17052 33368 17080 33467
rect 18708 33448 18736 33476
rect 18877 33473 18889 33507
rect 18923 33504 18935 33507
rect 21269 33507 21327 33513
rect 18923 33476 19564 33504
rect 18923 33473 18935 33476
rect 18877 33467 18935 33473
rect 19536 33448 19564 33476
rect 21269 33473 21281 33507
rect 21315 33473 21327 33507
rect 21269 33467 21327 33473
rect 22465 33507 22523 33513
rect 22465 33473 22477 33507
rect 22511 33504 22523 33507
rect 24026 33504 24032 33516
rect 22511 33476 24032 33504
rect 22511 33473 22523 33476
rect 22465 33467 22523 33473
rect 24026 33464 24032 33476
rect 24084 33464 24090 33516
rect 17586 33436 17592 33448
rect 17547 33408 17592 33436
rect 17586 33396 17592 33408
rect 17644 33396 17650 33448
rect 18690 33436 18696 33448
rect 18651 33408 18696 33436
rect 18690 33396 18696 33408
rect 18748 33396 18754 33448
rect 18785 33439 18843 33445
rect 18785 33405 18797 33439
rect 18831 33405 18843 33439
rect 18785 33399 18843 33405
rect 13924 33340 17080 33368
rect 17604 33368 17632 33396
rect 18800 33368 18828 33399
rect 18966 33396 18972 33448
rect 19024 33436 19030 33448
rect 19518 33436 19524 33448
rect 19024 33408 19069 33436
rect 19431 33408 19524 33436
rect 19024 33396 19030 33408
rect 19518 33396 19524 33408
rect 19576 33396 19582 33448
rect 20898 33396 20904 33448
rect 20956 33436 20962 33448
rect 20993 33439 21051 33445
rect 20993 33436 21005 33439
rect 20956 33408 21005 33436
rect 20956 33396 20962 33408
rect 20993 33405 21005 33408
rect 21039 33405 21051 33439
rect 20993 33399 21051 33405
rect 22189 33439 22247 33445
rect 22189 33405 22201 33439
rect 22235 33405 22247 33439
rect 23474 33436 23480 33448
rect 23435 33408 23480 33436
rect 22189 33399 22247 33405
rect 17604 33340 18828 33368
rect 22204 33368 22232 33399
rect 23474 33396 23480 33408
rect 23532 33396 23538 33448
rect 24412 33368 24440 33544
rect 25222 33532 25228 33544
rect 25280 33532 25286 33584
rect 30006 33532 30012 33584
rect 30064 33532 30070 33584
rect 30190 33532 30196 33584
rect 30248 33572 30254 33584
rect 30469 33575 30527 33581
rect 30469 33572 30481 33575
rect 30248 33544 30481 33572
rect 30248 33532 30254 33544
rect 30469 33541 30481 33544
rect 30515 33541 30527 33575
rect 30469 33535 30527 33541
rect 24489 33507 24547 33513
rect 24489 33473 24501 33507
rect 24535 33504 24547 33507
rect 24688 33504 24900 33510
rect 25038 33504 25044 33516
rect 24535 33482 25044 33504
rect 24535 33476 24716 33482
rect 24872 33476 25044 33482
rect 24535 33473 24547 33476
rect 24489 33467 24547 33473
rect 25038 33464 25044 33476
rect 25096 33464 25102 33516
rect 25590 33504 25596 33516
rect 25551 33476 25596 33504
rect 25590 33464 25596 33476
rect 25648 33464 25654 33516
rect 26970 33504 26976 33516
rect 26931 33476 26976 33504
rect 26970 33464 26976 33476
rect 27028 33464 27034 33516
rect 27890 33504 27896 33516
rect 27851 33476 27896 33504
rect 27890 33464 27896 33476
rect 27948 33464 27954 33516
rect 28077 33507 28135 33513
rect 28077 33473 28089 33507
rect 28123 33504 28135 33507
rect 28166 33504 28172 33516
rect 28123 33476 28172 33504
rect 28123 33473 28135 33476
rect 28077 33467 28135 33473
rect 28166 33464 28172 33476
rect 28224 33464 28230 33516
rect 32122 33504 32128 33516
rect 32083 33476 32128 33504
rect 32122 33464 32128 33476
rect 32180 33464 32186 33516
rect 32398 33464 32404 33516
rect 32456 33504 32462 33516
rect 33321 33507 33379 33513
rect 33321 33504 33333 33507
rect 32456 33476 33333 33504
rect 32456 33464 32462 33476
rect 33321 33473 33333 33476
rect 33367 33504 33379 33507
rect 34698 33504 34704 33516
rect 33367 33476 34704 33504
rect 33367 33473 33379 33476
rect 33321 33467 33379 33473
rect 34698 33464 34704 33476
rect 34756 33464 34762 33516
rect 36262 33464 36268 33516
rect 36320 33504 36326 33516
rect 36541 33507 36599 33513
rect 36541 33504 36553 33507
rect 36320 33476 36553 33504
rect 36320 33464 36326 33476
rect 36541 33473 36553 33476
rect 36587 33473 36599 33507
rect 36541 33467 36599 33473
rect 37461 33507 37519 33513
rect 37461 33473 37473 33507
rect 37507 33473 37519 33507
rect 38102 33504 38108 33516
rect 38063 33476 38108 33504
rect 37461 33467 37519 33473
rect 24578 33436 24584 33448
rect 24539 33408 24584 33436
rect 24578 33396 24584 33408
rect 24636 33396 24642 33448
rect 24673 33439 24731 33445
rect 24673 33436 24685 33439
rect 24672 33405 24685 33436
rect 24719 33405 24731 33439
rect 24672 33399 24731 33405
rect 24768 33439 24826 33445
rect 24768 33405 24780 33439
rect 24814 33405 24826 33439
rect 24768 33399 24826 33405
rect 22204 33340 24440 33368
rect 16758 33300 16764 33312
rect 11348 33272 16764 33300
rect 16758 33260 16764 33272
rect 16816 33260 16822 33312
rect 17773 33303 17831 33309
rect 17773 33269 17785 33303
rect 17819 33300 17831 33303
rect 18598 33300 18604 33312
rect 17819 33272 18604 33300
rect 17819 33269 17831 33272
rect 17773 33263 17831 33269
rect 18598 33260 18604 33272
rect 18656 33260 18662 33312
rect 22373 33303 22431 33309
rect 22373 33269 22385 33303
rect 22419 33300 22431 33303
rect 23566 33300 23572 33312
rect 22419 33272 23572 33300
rect 22419 33269 22431 33272
rect 22373 33263 22431 33269
rect 23566 33260 23572 33272
rect 23624 33260 23630 33312
rect 24394 33260 24400 33312
rect 24452 33300 24458 33312
rect 24672 33300 24700 33399
rect 24452 33272 24700 33300
rect 24780 33300 24808 33399
rect 24854 33396 24860 33448
rect 24912 33436 24918 33448
rect 25406 33436 25412 33448
rect 24912 33408 25412 33436
rect 24912 33396 24918 33408
rect 25406 33396 25412 33408
rect 25464 33396 25470 33448
rect 27798 33436 27804 33448
rect 27759 33408 27804 33436
rect 27798 33396 27804 33408
rect 27856 33396 27862 33448
rect 27982 33396 27988 33448
rect 28040 33436 28046 33448
rect 30745 33439 30803 33445
rect 28040 33408 28085 33436
rect 28040 33396 28046 33408
rect 30745 33405 30757 33439
rect 30791 33436 30803 33439
rect 30926 33436 30932 33448
rect 30791 33408 30932 33436
rect 30791 33405 30803 33408
rect 30745 33399 30803 33405
rect 30926 33396 30932 33408
rect 30984 33396 30990 33448
rect 31018 33396 31024 33448
rect 31076 33436 31082 33448
rect 37476 33436 37504 33467
rect 38102 33464 38108 33476
rect 38160 33464 38166 33516
rect 37550 33436 37556 33448
rect 31076 33408 37556 33436
rect 31076 33396 31082 33408
rect 37550 33396 37556 33408
rect 37608 33396 37614 33448
rect 24946 33300 24952 33312
rect 24780 33272 24952 33300
rect 24452 33260 24458 33272
rect 24946 33260 24952 33272
rect 25004 33260 25010 33312
rect 27062 33300 27068 33312
rect 27023 33272 27068 33300
rect 27062 33260 27068 33272
rect 27120 33260 27126 33312
rect 28994 33300 29000 33312
rect 28955 33272 29000 33300
rect 28994 33260 29000 33272
rect 29052 33260 29058 33312
rect 30834 33260 30840 33312
rect 30892 33300 30898 33312
rect 31754 33300 31760 33312
rect 30892 33272 31760 33300
rect 30892 33260 30898 33272
rect 31754 33260 31760 33272
rect 31812 33260 31818 33312
rect 32030 33260 32036 33312
rect 32088 33300 32094 33312
rect 32309 33303 32367 33309
rect 32309 33300 32321 33303
rect 32088 33272 32321 33300
rect 32088 33260 32094 33272
rect 32309 33269 32321 33272
rect 32355 33300 32367 33303
rect 32950 33300 32956 33312
rect 32355 33272 32956 33300
rect 32355 33269 32367 33272
rect 32309 33263 32367 33269
rect 32950 33260 32956 33272
rect 33008 33260 33014 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 8941 33099 8999 33105
rect 8941 33065 8953 33099
rect 8987 33096 8999 33099
rect 10318 33096 10324 33108
rect 8987 33068 10324 33096
rect 8987 33065 8999 33068
rect 8941 33059 8999 33065
rect 10318 33056 10324 33068
rect 10376 33056 10382 33108
rect 11238 33056 11244 33108
rect 11296 33096 11302 33108
rect 12805 33099 12863 33105
rect 11296 33068 12434 33096
rect 11296 33056 11302 33068
rect 10870 32988 10876 33040
rect 10928 33028 10934 33040
rect 10928 33000 12204 33028
rect 10928 32988 10934 33000
rect 7561 32963 7619 32969
rect 7561 32929 7573 32963
rect 7607 32929 7619 32963
rect 7561 32923 7619 32929
rect 5810 32892 5816 32904
rect 5771 32864 5816 32892
rect 5810 32852 5816 32864
rect 5868 32852 5874 32904
rect 4706 32784 4712 32836
rect 4764 32824 4770 32836
rect 5261 32827 5319 32833
rect 5261 32824 5273 32827
rect 4764 32796 5273 32824
rect 4764 32784 4770 32796
rect 5261 32793 5273 32796
rect 5307 32793 5319 32827
rect 7576 32824 7604 32923
rect 8478 32920 8484 32972
rect 8536 32960 8542 32972
rect 10689 32963 10747 32969
rect 10689 32960 10701 32963
rect 8536 32932 10701 32960
rect 8536 32920 8542 32932
rect 10689 32929 10701 32932
rect 10735 32960 10747 32963
rect 11514 32960 11520 32972
rect 10735 32932 11520 32960
rect 10735 32929 10747 32932
rect 10689 32923 10747 32929
rect 11514 32920 11520 32932
rect 11572 32920 11578 32972
rect 7742 32892 7748 32904
rect 7703 32864 7748 32892
rect 7742 32852 7748 32864
rect 7800 32852 7806 32904
rect 7834 32852 7840 32904
rect 7892 32892 7898 32904
rect 11333 32895 11391 32901
rect 7892 32864 7937 32892
rect 7892 32852 7898 32864
rect 11333 32861 11345 32895
rect 11379 32861 11391 32895
rect 11333 32855 11391 32861
rect 11425 32895 11483 32901
rect 11425 32861 11437 32895
rect 11471 32861 11483 32895
rect 11606 32892 11612 32904
rect 11567 32864 11612 32892
rect 11425 32855 11483 32861
rect 7576 32796 9076 32824
rect 5261 32787 5319 32793
rect 7374 32716 7380 32768
rect 7432 32756 7438 32768
rect 7561 32759 7619 32765
rect 7561 32756 7573 32759
rect 7432 32728 7573 32756
rect 7432 32716 7438 32728
rect 7561 32725 7573 32728
rect 7607 32725 7619 32759
rect 9048 32756 9076 32796
rect 9122 32784 9128 32836
rect 9180 32824 9186 32836
rect 10410 32824 10416 32836
rect 9180 32796 9246 32824
rect 10371 32796 10416 32824
rect 9180 32784 9186 32796
rect 10410 32784 10416 32796
rect 10468 32784 10474 32836
rect 9766 32756 9772 32768
rect 9048 32728 9772 32756
rect 7561 32719 7619 32725
rect 9766 32716 9772 32728
rect 9824 32716 9830 32768
rect 10042 32716 10048 32768
rect 10100 32756 10106 32768
rect 11149 32759 11207 32765
rect 11149 32756 11161 32759
rect 10100 32728 11161 32756
rect 10100 32716 10106 32728
rect 11149 32725 11161 32728
rect 11195 32725 11207 32759
rect 11348 32756 11376 32855
rect 11440 32824 11468 32855
rect 11606 32852 11612 32864
rect 11664 32852 11670 32904
rect 11701 32895 11759 32901
rect 11701 32861 11713 32895
rect 11747 32892 11759 32895
rect 11882 32892 11888 32904
rect 11747 32864 11888 32892
rect 11747 32861 11759 32864
rect 11701 32855 11759 32861
rect 11882 32852 11888 32864
rect 11940 32852 11946 32904
rect 12176 32901 12204 33000
rect 12406 32960 12434 33068
rect 12805 33065 12817 33099
rect 12851 33096 12863 33099
rect 12894 33096 12900 33108
rect 12851 33068 12900 33096
rect 12851 33065 12863 33068
rect 12805 33059 12863 33065
rect 12894 33056 12900 33068
rect 12952 33056 12958 33108
rect 14642 33056 14648 33108
rect 14700 33096 14706 33108
rect 14829 33099 14887 33105
rect 14829 33096 14841 33099
rect 14700 33068 14841 33096
rect 14700 33056 14706 33068
rect 14829 33065 14841 33068
rect 14875 33096 14887 33099
rect 18414 33096 18420 33108
rect 14875 33068 16804 33096
rect 18375 33068 18420 33096
rect 14875 33065 14887 33068
rect 14829 33059 14887 33065
rect 14274 33028 14280 33040
rect 13464 33000 14280 33028
rect 13464 32969 13492 33000
rect 14274 32988 14280 33000
rect 14332 32988 14338 33040
rect 16776 33028 16804 33068
rect 18414 33056 18420 33068
rect 18472 33056 18478 33108
rect 20714 33096 20720 33108
rect 20675 33068 20720 33096
rect 20714 33056 20720 33068
rect 20772 33056 20778 33108
rect 22646 33056 22652 33108
rect 22704 33096 22710 33108
rect 22741 33099 22799 33105
rect 22741 33096 22753 33099
rect 22704 33068 22753 33096
rect 22704 33056 22710 33068
rect 22741 33065 22753 33068
rect 22787 33065 22799 33099
rect 22741 33059 22799 33065
rect 23569 33099 23627 33105
rect 23569 33065 23581 33099
rect 23615 33096 23627 33099
rect 24578 33096 24584 33108
rect 23615 33068 24584 33096
rect 23615 33065 23627 33068
rect 23569 33059 23627 33065
rect 24578 33056 24584 33068
rect 24636 33056 24642 33108
rect 24673 33099 24731 33105
rect 24673 33065 24685 33099
rect 24719 33065 24731 33099
rect 27801 33099 27859 33105
rect 24673 33059 24731 33065
rect 24780 33068 27384 33096
rect 19797 33031 19855 33037
rect 16776 33000 19656 33028
rect 12989 32963 13047 32969
rect 12989 32960 13001 32963
rect 12406 32932 13001 32960
rect 12989 32929 13001 32932
rect 13035 32929 13047 32963
rect 12989 32923 13047 32929
rect 13449 32963 13507 32969
rect 13449 32929 13461 32963
rect 13495 32929 13507 32963
rect 13449 32923 13507 32929
rect 15378 32920 15384 32972
rect 15436 32960 15442 32972
rect 15473 32963 15531 32969
rect 15473 32960 15485 32963
rect 15436 32932 15485 32960
rect 15436 32920 15442 32932
rect 15473 32929 15485 32932
rect 15519 32929 15531 32963
rect 15473 32923 15531 32929
rect 18230 32920 18236 32972
rect 18288 32960 18294 32972
rect 18325 32963 18383 32969
rect 18325 32960 18337 32963
rect 18288 32932 18337 32960
rect 18288 32920 18294 32932
rect 18325 32929 18337 32932
rect 18371 32929 18383 32963
rect 18325 32923 18383 32929
rect 12161 32895 12219 32901
rect 12161 32861 12173 32895
rect 12207 32861 12219 32895
rect 13078 32892 13084 32904
rect 13039 32864 13084 32892
rect 12161 32855 12219 32861
rect 13078 32852 13084 32864
rect 13136 32852 13142 32904
rect 13998 32852 14004 32904
rect 14056 32892 14062 32904
rect 14277 32895 14335 32901
rect 14277 32892 14289 32895
rect 14056 32864 14289 32892
rect 14056 32852 14062 32864
rect 14277 32861 14289 32864
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 14921 32895 14979 32901
rect 14921 32861 14933 32895
rect 14967 32892 14979 32895
rect 15286 32892 15292 32904
rect 14967 32864 15292 32892
rect 14967 32861 14979 32864
rect 14921 32855 14979 32861
rect 15286 32852 15292 32864
rect 15344 32852 15350 32904
rect 18414 32892 18420 32904
rect 16882 32864 18420 32892
rect 18414 32852 18420 32864
rect 18472 32852 18478 32904
rect 18509 32895 18567 32901
rect 18509 32861 18521 32895
rect 18555 32892 18567 32895
rect 18966 32892 18972 32904
rect 18555 32864 18972 32892
rect 18555 32861 18567 32864
rect 18509 32855 18567 32861
rect 18966 32852 18972 32864
rect 19024 32852 19030 32904
rect 19150 32852 19156 32904
rect 19208 32892 19214 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 19208 32864 19257 32892
rect 19208 32852 19214 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19518 32892 19524 32904
rect 19479 32864 19524 32892
rect 19245 32855 19303 32861
rect 19518 32852 19524 32864
rect 19576 32852 19582 32904
rect 19628 32901 19656 33000
rect 19797 32997 19809 33031
rect 19843 33028 19855 33031
rect 20898 33028 20904 33040
rect 19843 33000 20904 33028
rect 19843 32997 19855 33000
rect 19797 32991 19855 32997
rect 20898 32988 20904 33000
rect 20956 32988 20962 33040
rect 24394 32988 24400 33040
rect 24452 33028 24458 33040
rect 24687 33028 24715 33059
rect 24452 33000 24715 33028
rect 24452 32988 24458 33000
rect 24780 32960 24808 33068
rect 27356 33028 27384 33068
rect 27801 33065 27813 33099
rect 27847 33096 27859 33099
rect 28166 33096 28172 33108
rect 27847 33068 28172 33096
rect 27847 33065 27859 33068
rect 27801 33059 27859 33065
rect 28166 33056 28172 33068
rect 28224 33056 28230 33108
rect 28534 33056 28540 33108
rect 28592 33096 28598 33108
rect 28629 33099 28687 33105
rect 28629 33096 28641 33099
rect 28592 33068 28641 33096
rect 28592 33056 28598 33068
rect 28629 33065 28641 33068
rect 28675 33065 28687 33099
rect 30190 33096 30196 33108
rect 30151 33068 30196 33096
rect 28629 33059 28687 33065
rect 30190 33056 30196 33068
rect 30248 33056 30254 33108
rect 30650 33096 30656 33108
rect 30611 33068 30656 33096
rect 30650 33056 30656 33068
rect 30708 33056 30714 33108
rect 30742 33056 30748 33108
rect 30800 33096 30806 33108
rect 31570 33096 31576 33108
rect 30800 33068 31576 33096
rect 30800 33056 30806 33068
rect 31018 33028 31024 33040
rect 27356 33000 31024 33028
rect 31018 32988 31024 33000
rect 31076 32988 31082 33040
rect 26050 32960 26056 32972
rect 22066 32932 24808 32960
rect 26011 32932 26056 32960
rect 19613 32895 19671 32901
rect 19613 32861 19625 32895
rect 19659 32892 19671 32895
rect 20070 32892 20076 32904
rect 19659 32864 20076 32892
rect 19659 32861 19671 32864
rect 19613 32855 19671 32861
rect 20070 32852 20076 32864
rect 20128 32852 20134 32904
rect 20806 32892 20812 32904
rect 20767 32864 20812 32892
rect 20806 32852 20812 32864
rect 20864 32852 20870 32904
rect 21361 32895 21419 32901
rect 21361 32861 21373 32895
rect 21407 32892 21419 32895
rect 21450 32892 21456 32904
rect 21407 32864 21456 32892
rect 21407 32861 21419 32864
rect 21361 32855 21419 32861
rect 21450 32852 21456 32864
rect 21508 32852 21514 32904
rect 12253 32827 12311 32833
rect 12253 32824 12265 32827
rect 11440 32796 12265 32824
rect 12253 32793 12265 32796
rect 12299 32793 12311 32827
rect 12253 32787 12311 32793
rect 13357 32827 13415 32833
rect 13357 32793 13369 32827
rect 13403 32824 13415 32827
rect 14642 32824 14648 32836
rect 13403 32796 14648 32824
rect 13403 32793 13415 32796
rect 13357 32787 13415 32793
rect 14642 32784 14648 32796
rect 14700 32784 14706 32836
rect 15194 32784 15200 32836
rect 15252 32824 15258 32836
rect 15749 32827 15807 32833
rect 15749 32824 15761 32827
rect 15252 32796 15761 32824
rect 15252 32784 15258 32796
rect 15749 32793 15761 32796
rect 15795 32793 15807 32827
rect 15749 32787 15807 32793
rect 17034 32784 17040 32836
rect 17092 32824 17098 32836
rect 18233 32827 18291 32833
rect 18233 32824 18245 32827
rect 17092 32796 18245 32824
rect 17092 32784 17098 32796
rect 18233 32793 18245 32796
rect 18279 32793 18291 32827
rect 18233 32787 18291 32793
rect 18598 32784 18604 32836
rect 18656 32824 18662 32836
rect 19429 32827 19487 32833
rect 19429 32824 19441 32827
rect 18656 32796 19441 32824
rect 18656 32784 18662 32796
rect 19429 32793 19441 32796
rect 19475 32793 19487 32827
rect 21726 32824 21732 32836
rect 21687 32796 21732 32824
rect 19429 32787 19487 32793
rect 21726 32784 21732 32796
rect 21784 32824 21790 32836
rect 22066 32824 22094 32932
rect 26050 32920 26056 32932
rect 26108 32920 26114 32972
rect 26326 32960 26332 32972
rect 26287 32932 26332 32960
rect 26326 32920 26332 32932
rect 26384 32920 26390 32972
rect 26418 32920 26424 32972
rect 26476 32960 26482 32972
rect 26476 32932 27844 32960
rect 26476 32920 26482 32932
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32892 22707 32895
rect 23382 32892 23388 32904
rect 22695 32864 23388 32892
rect 22695 32861 22707 32864
rect 22649 32855 22707 32861
rect 23382 32852 23388 32864
rect 23440 32852 23446 32904
rect 23474 32852 23480 32904
rect 23532 32852 23538 32904
rect 24486 32852 24492 32904
rect 24544 32892 24550 32904
rect 25409 32895 25467 32901
rect 25409 32892 25421 32895
rect 24544 32864 25421 32892
rect 24544 32852 24550 32864
rect 25409 32861 25421 32864
rect 25455 32861 25467 32895
rect 27816 32892 27844 32932
rect 27890 32920 27896 32972
rect 27948 32960 27954 32972
rect 30466 32960 30472 32972
rect 27948 32932 30472 32960
rect 27948 32920 27954 32932
rect 30466 32920 30472 32932
rect 30524 32920 30530 32972
rect 28534 32892 28540 32904
rect 27816 32864 28540 32892
rect 25409 32855 25467 32861
rect 28534 32852 28540 32864
rect 28592 32852 28598 32904
rect 28629 32895 28687 32901
rect 28629 32861 28641 32895
rect 28675 32861 28687 32895
rect 28629 32855 28687 32861
rect 21784 32796 22094 32824
rect 23492 32824 23520 32852
rect 23753 32827 23811 32833
rect 23753 32824 23765 32827
rect 23492 32796 23765 32824
rect 21784 32784 21790 32796
rect 23753 32793 23765 32796
rect 23799 32824 23811 32827
rect 24302 32824 24308 32836
rect 23799 32796 24308 32824
rect 23799 32793 23811 32796
rect 23753 32787 23811 32793
rect 24302 32784 24308 32796
rect 24360 32784 24366 32836
rect 24857 32827 24915 32833
rect 24857 32793 24869 32827
rect 24903 32824 24915 32827
rect 25038 32824 25044 32836
rect 24903 32796 25044 32824
rect 24903 32793 24915 32796
rect 24857 32787 24915 32793
rect 25038 32784 25044 32796
rect 25096 32784 25102 32836
rect 25424 32796 26740 32824
rect 11790 32756 11796 32768
rect 11348 32728 11796 32756
rect 11149 32719 11207 32725
rect 11790 32716 11796 32728
rect 11848 32716 11854 32768
rect 14182 32756 14188 32768
rect 14143 32728 14188 32756
rect 14182 32716 14188 32728
rect 14240 32716 14246 32768
rect 16482 32716 16488 32768
rect 16540 32756 16546 32768
rect 17221 32759 17279 32765
rect 17221 32756 17233 32759
rect 16540 32728 17233 32756
rect 16540 32716 16546 32728
rect 17221 32725 17233 32728
rect 17267 32725 17279 32759
rect 17221 32719 17279 32725
rect 18322 32716 18328 32768
rect 18380 32756 18386 32768
rect 18693 32759 18751 32765
rect 18693 32756 18705 32759
rect 18380 32728 18705 32756
rect 18380 32716 18386 32728
rect 18693 32725 18705 32728
rect 18739 32725 18751 32759
rect 18693 32719 18751 32725
rect 22922 32716 22928 32768
rect 22980 32756 22986 32768
rect 23566 32765 23572 32768
rect 23385 32759 23443 32765
rect 23385 32756 23397 32759
rect 22980 32728 23397 32756
rect 22980 32716 22986 32728
rect 23385 32725 23397 32728
rect 23431 32725 23443 32759
rect 23385 32719 23443 32725
rect 23553 32759 23572 32765
rect 23553 32725 23565 32759
rect 23624 32756 23630 32768
rect 24210 32756 24216 32768
rect 23624 32728 24216 32756
rect 23553 32719 23572 32725
rect 23566 32716 23572 32719
rect 23624 32716 23630 32728
rect 24210 32716 24216 32728
rect 24268 32756 24274 32768
rect 24489 32759 24547 32765
rect 24489 32756 24501 32759
rect 24268 32728 24501 32756
rect 24268 32716 24274 32728
rect 24489 32725 24501 32728
rect 24535 32725 24547 32759
rect 24489 32719 24547 32725
rect 24657 32759 24715 32765
rect 24657 32725 24669 32759
rect 24703 32756 24715 32759
rect 24946 32756 24952 32768
rect 24703 32728 24952 32756
rect 24703 32725 24715 32728
rect 24657 32719 24715 32725
rect 24946 32716 24952 32728
rect 25004 32756 25010 32768
rect 25424 32756 25452 32796
rect 25004 32728 25452 32756
rect 25004 32716 25010 32728
rect 25498 32716 25504 32768
rect 25556 32756 25562 32768
rect 26418 32756 26424 32768
rect 25556 32728 26424 32756
rect 25556 32716 25562 32728
rect 26418 32716 26424 32728
rect 26476 32716 26482 32768
rect 26712 32756 26740 32796
rect 27062 32784 27068 32836
rect 27120 32784 27126 32836
rect 28644 32824 28672 32855
rect 28718 32852 28724 32904
rect 28776 32892 28782 32904
rect 28994 32892 29000 32904
rect 28776 32864 29000 32892
rect 28776 32852 28782 32864
rect 28994 32852 29000 32864
rect 29052 32892 29058 32904
rect 29822 32892 29828 32904
rect 29052 32864 29828 32892
rect 29052 32852 29058 32864
rect 29822 32852 29828 32864
rect 29880 32892 29886 32904
rect 29917 32895 29975 32901
rect 29917 32892 29929 32895
rect 29880 32864 29929 32892
rect 29880 32852 29886 32864
rect 29917 32861 29929 32864
rect 29963 32861 29975 32895
rect 29917 32855 29975 32861
rect 30009 32895 30067 32901
rect 30009 32861 30021 32895
rect 30055 32892 30067 32895
rect 30098 32892 30104 32904
rect 30055 32864 30104 32892
rect 30055 32861 30067 32864
rect 30009 32855 30067 32861
rect 30098 32852 30104 32864
rect 30156 32852 30162 32904
rect 30834 32892 30840 32904
rect 30795 32864 30840 32892
rect 30834 32852 30840 32864
rect 30892 32852 30898 32904
rect 31174 32901 31202 33068
rect 31570 33056 31576 33068
rect 31628 33056 31634 33108
rect 31754 33096 31760 33108
rect 31715 33068 31760 33096
rect 31754 33056 31760 33068
rect 31812 33056 31818 33108
rect 31846 33056 31852 33108
rect 31904 33096 31910 33108
rect 33594 33096 33600 33108
rect 31904 33068 33600 33096
rect 31904 33056 31910 33068
rect 33594 33056 33600 33068
rect 33652 33056 33658 33108
rect 31938 32960 31944 32972
rect 31899 32932 31944 32960
rect 31938 32920 31944 32932
rect 31996 32920 32002 32972
rect 32140 32969 32352 32976
rect 32125 32963 32352 32969
rect 32125 32929 32137 32963
rect 32171 32960 32352 32963
rect 32490 32960 32496 32972
rect 32171 32948 32496 32960
rect 32171 32929 32183 32948
rect 32324 32932 32496 32948
rect 32125 32923 32183 32929
rect 32490 32920 32496 32932
rect 32548 32960 32554 32972
rect 32548 32932 34008 32960
rect 32548 32920 32554 32932
rect 31021 32895 31079 32901
rect 31021 32882 31033 32895
rect 31067 32882 31079 32895
rect 31159 32895 31217 32901
rect 30929 32827 30987 32833
rect 31018 32830 31024 32882
rect 31076 32830 31082 32882
rect 31159 32861 31171 32895
rect 31205 32861 31217 32895
rect 31159 32855 31217 32861
rect 31294 32852 31300 32904
rect 31352 32892 31358 32904
rect 32030 32892 32036 32904
rect 31352 32864 31397 32892
rect 31991 32864 32036 32892
rect 31352 32852 31358 32864
rect 32030 32852 32036 32864
rect 32088 32852 32094 32904
rect 32232 32901 32444 32902
rect 32217 32895 32444 32901
rect 32217 32861 32229 32895
rect 32263 32874 32444 32895
rect 32766 32892 32772 32904
rect 32263 32861 32275 32874
rect 32217 32855 32275 32861
rect 30929 32824 30941 32827
rect 28644 32796 30941 32824
rect 30929 32793 30941 32796
rect 30975 32793 30987 32827
rect 30929 32787 30987 32793
rect 28442 32756 28448 32768
rect 26712 32728 28448 32756
rect 28442 32716 28448 32728
rect 28500 32716 28506 32768
rect 28997 32759 29055 32765
rect 28997 32725 29009 32759
rect 29043 32756 29055 32759
rect 29549 32759 29607 32765
rect 29549 32756 29561 32759
rect 29043 32728 29561 32756
rect 29043 32725 29055 32728
rect 28997 32719 29055 32725
rect 29549 32725 29561 32728
rect 29595 32725 29607 32759
rect 30944 32756 30972 32787
rect 31570 32784 31576 32836
rect 31628 32824 31634 32836
rect 32416 32824 32444 32874
rect 32727 32864 32772 32892
rect 32766 32852 32772 32864
rect 32824 32852 32830 32904
rect 33980 32901 34008 32932
rect 33965 32895 34023 32901
rect 33965 32861 33977 32895
rect 34011 32861 34023 32895
rect 34698 32892 34704 32904
rect 34659 32864 34704 32892
rect 33965 32855 34023 32861
rect 34698 32852 34704 32864
rect 34756 32852 34762 32904
rect 36262 32892 36268 32904
rect 36223 32864 36268 32892
rect 36262 32852 36268 32864
rect 36320 32852 36326 32904
rect 31628 32796 32444 32824
rect 31628 32784 31634 32796
rect 32950 32784 32956 32836
rect 33008 32824 33014 32836
rect 33008 32796 33053 32824
rect 33008 32784 33014 32796
rect 33686 32784 33692 32836
rect 33744 32824 33750 32836
rect 33781 32827 33839 32833
rect 33781 32824 33793 32827
rect 33744 32796 33793 32824
rect 33744 32784 33750 32796
rect 33781 32793 33793 32796
rect 33827 32793 33839 32827
rect 33781 32787 33839 32793
rect 36449 32827 36507 32833
rect 36449 32793 36461 32827
rect 36495 32824 36507 32827
rect 37642 32824 37648 32836
rect 36495 32796 37648 32824
rect 36495 32793 36507 32796
rect 36449 32787 36507 32793
rect 37642 32784 37648 32796
rect 37700 32784 37706 32836
rect 38102 32824 38108 32836
rect 38063 32796 38108 32824
rect 38102 32784 38108 32796
rect 38160 32784 38166 32836
rect 31754 32756 31760 32768
rect 30944 32728 31760 32756
rect 29549 32719 29607 32725
rect 31754 32716 31760 32728
rect 31812 32716 31818 32768
rect 32398 32716 32404 32768
rect 32456 32756 32462 32768
rect 33137 32759 33195 32765
rect 33137 32756 33149 32759
rect 32456 32728 33149 32756
rect 32456 32716 32462 32728
rect 33137 32725 33149 32728
rect 33183 32725 33195 32759
rect 33137 32719 33195 32725
rect 34054 32716 34060 32768
rect 34112 32756 34118 32768
rect 34149 32759 34207 32765
rect 34149 32756 34161 32759
rect 34112 32728 34161 32756
rect 34112 32716 34118 32728
rect 34149 32725 34161 32728
rect 34195 32725 34207 32759
rect 34790 32756 34796 32768
rect 34751 32728 34796 32756
rect 34149 32719 34207 32725
rect 34790 32716 34796 32728
rect 34848 32716 34854 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 8478 32552 8484 32564
rect 7484 32524 8484 32552
rect 6730 32484 6736 32496
rect 5828 32456 6736 32484
rect 5828 32425 5856 32456
rect 6730 32444 6736 32456
rect 6788 32444 6794 32496
rect 5813 32419 5871 32425
rect 5813 32385 5825 32419
rect 5859 32385 5871 32419
rect 6822 32416 6828 32428
rect 6783 32388 6828 32416
rect 5813 32379 5871 32385
rect 6822 32376 6828 32388
rect 6880 32376 6886 32428
rect 7006 32416 7012 32428
rect 6967 32388 7012 32416
rect 7006 32376 7012 32388
rect 7064 32376 7070 32428
rect 6546 32308 6552 32360
rect 6604 32348 6610 32360
rect 7484 32357 7512 32524
rect 8478 32512 8484 32524
rect 8536 32512 8542 32564
rect 10244 32524 10364 32552
rect 8386 32444 8392 32496
rect 8444 32444 8450 32496
rect 10244 32493 10272 32524
rect 10229 32487 10287 32493
rect 10229 32453 10241 32487
rect 10275 32453 10287 32487
rect 10336 32484 10364 32524
rect 10410 32512 10416 32564
rect 10468 32552 10474 32564
rect 11517 32555 11575 32561
rect 11517 32552 11529 32555
rect 10468 32524 11529 32552
rect 10468 32512 10474 32524
rect 11517 32521 11529 32524
rect 11563 32521 11575 32555
rect 11517 32515 11575 32521
rect 12802 32512 12808 32564
rect 12860 32552 12866 32564
rect 13078 32552 13084 32564
rect 12860 32524 13084 32552
rect 12860 32512 12866 32524
rect 13078 32512 13084 32524
rect 13136 32512 13142 32564
rect 15194 32552 15200 32564
rect 15155 32524 15200 32552
rect 15194 32512 15200 32524
rect 15252 32512 15258 32564
rect 15378 32512 15384 32564
rect 15436 32552 15442 32564
rect 17957 32555 18015 32561
rect 17957 32552 17969 32555
rect 15436 32524 17969 32552
rect 15436 32512 15442 32524
rect 17957 32521 17969 32524
rect 18003 32552 18015 32555
rect 19242 32552 19248 32564
rect 18003 32524 19248 32552
rect 18003 32521 18015 32524
rect 17957 32515 18015 32521
rect 19242 32512 19248 32524
rect 19300 32552 19306 32564
rect 20990 32552 20996 32564
rect 19300 32524 20996 32552
rect 19300 32512 19306 32524
rect 20990 32512 20996 32524
rect 21048 32512 21054 32564
rect 21269 32555 21327 32561
rect 21269 32521 21281 32555
rect 21315 32552 21327 32555
rect 25317 32555 25375 32561
rect 21315 32524 22140 32552
rect 21315 32521 21327 32524
rect 21269 32515 21327 32521
rect 11054 32484 11060 32496
rect 10336 32456 11060 32484
rect 10229 32447 10287 32453
rect 11054 32444 11060 32456
rect 11112 32444 11118 32496
rect 11885 32487 11943 32493
rect 11885 32453 11897 32487
rect 11931 32484 11943 32487
rect 12986 32484 12992 32496
rect 11931 32456 12992 32484
rect 11931 32453 11943 32456
rect 11885 32447 11943 32453
rect 12986 32444 12992 32456
rect 13044 32444 13050 32496
rect 13173 32487 13231 32493
rect 13173 32453 13185 32487
rect 13219 32484 13231 32487
rect 13817 32487 13875 32493
rect 13817 32484 13829 32487
rect 13219 32456 13829 32484
rect 13219 32453 13231 32456
rect 13173 32447 13231 32453
rect 13817 32453 13829 32456
rect 13863 32484 13875 32487
rect 14553 32487 14611 32493
rect 14553 32484 14565 32487
rect 13863 32456 14565 32484
rect 13863 32453 13875 32456
rect 13817 32447 13875 32453
rect 14553 32453 14565 32456
rect 14599 32484 14611 32487
rect 15286 32484 15292 32496
rect 14599 32456 15292 32484
rect 14599 32453 14611 32456
rect 14553 32447 14611 32453
rect 15286 32444 15292 32456
rect 15344 32444 15350 32496
rect 15470 32484 15476 32496
rect 15431 32456 15476 32484
rect 15470 32444 15476 32456
rect 15528 32484 15534 32496
rect 16482 32484 16488 32496
rect 15528 32456 16488 32484
rect 15528 32444 15534 32456
rect 16482 32444 16488 32456
rect 16540 32484 16546 32496
rect 19061 32487 19119 32493
rect 16540 32456 17080 32484
rect 16540 32444 16546 32456
rect 9953 32419 10011 32425
rect 9953 32385 9965 32419
rect 9999 32416 10011 32419
rect 10042 32416 10048 32428
rect 9999 32388 10048 32416
rect 9999 32385 10011 32388
rect 9953 32379 10011 32385
rect 10042 32376 10048 32388
rect 10100 32376 10106 32428
rect 10410 32376 10416 32428
rect 10468 32416 10474 32428
rect 10781 32419 10839 32425
rect 10781 32416 10793 32419
rect 10468 32388 10793 32416
rect 10468 32376 10474 32388
rect 10781 32385 10793 32388
rect 10827 32385 10839 32419
rect 11698 32416 11704 32428
rect 11659 32388 11704 32416
rect 10781 32379 10839 32385
rect 11698 32376 11704 32388
rect 11756 32376 11762 32428
rect 11790 32376 11796 32428
rect 11848 32416 11854 32428
rect 12023 32419 12081 32425
rect 11848 32388 11893 32416
rect 11848 32376 11854 32388
rect 12023 32385 12035 32419
rect 12069 32416 12081 32419
rect 12250 32416 12256 32428
rect 12069 32388 12256 32416
rect 12069 32385 12081 32388
rect 12023 32379 12081 32385
rect 12250 32376 12256 32388
rect 12308 32416 12314 32428
rect 14001 32419 14059 32425
rect 14001 32416 14013 32419
rect 12308 32388 14013 32416
rect 12308 32376 12314 32388
rect 14001 32385 14013 32388
rect 14047 32416 14059 32419
rect 15378 32416 15384 32428
rect 14047 32388 15384 32416
rect 14047 32385 14059 32388
rect 14001 32379 14059 32385
rect 15378 32376 15384 32388
rect 15436 32376 15442 32428
rect 15562 32416 15568 32428
rect 15523 32388 15568 32416
rect 15562 32376 15568 32388
rect 15620 32376 15626 32428
rect 17052 32425 17080 32456
rect 19061 32453 19073 32487
rect 19107 32484 19119 32487
rect 19426 32484 19432 32496
rect 19107 32456 19432 32484
rect 19107 32453 19119 32456
rect 19061 32447 19119 32453
rect 19426 32444 19432 32456
rect 19484 32444 19490 32496
rect 21008 32484 21036 32512
rect 22112 32493 22140 32524
rect 25317 32521 25329 32555
rect 25363 32552 25375 32555
rect 25958 32552 25964 32564
rect 25363 32524 25964 32552
rect 25363 32521 25375 32524
rect 25317 32515 25375 32521
rect 25958 32512 25964 32524
rect 26016 32512 26022 32564
rect 26237 32555 26295 32561
rect 26237 32521 26249 32555
rect 26283 32552 26295 32555
rect 26970 32552 26976 32564
rect 26283 32524 26976 32552
rect 26283 32521 26295 32524
rect 26237 32515 26295 32521
rect 26970 32512 26976 32524
rect 27028 32512 27034 32564
rect 27798 32561 27804 32564
rect 27785 32555 27804 32561
rect 27785 32552 27797 32555
rect 27711 32524 27797 32552
rect 27785 32521 27797 32524
rect 27856 32552 27862 32564
rect 28613 32555 28671 32561
rect 28613 32552 28625 32555
rect 27856 32524 28625 32552
rect 27785 32515 27804 32521
rect 27798 32512 27804 32515
rect 27856 32512 27862 32524
rect 28613 32521 28625 32524
rect 28659 32552 28671 32555
rect 28902 32552 28908 32564
rect 28659 32524 28908 32552
rect 28659 32521 28671 32524
rect 28613 32515 28671 32521
rect 28902 32512 28908 32524
rect 28960 32512 28966 32564
rect 30098 32552 30104 32564
rect 30059 32524 30104 32552
rect 30098 32512 30104 32524
rect 30156 32512 30162 32564
rect 30650 32512 30656 32564
rect 30708 32552 30714 32564
rect 31021 32555 31079 32561
rect 31021 32552 31033 32555
rect 30708 32524 31033 32552
rect 30708 32512 30714 32524
rect 31021 32521 31033 32524
rect 31067 32521 31079 32555
rect 31021 32515 31079 32521
rect 31205 32555 31263 32561
rect 31205 32521 31217 32555
rect 31251 32552 31263 32555
rect 32030 32552 32036 32564
rect 31251 32524 32036 32552
rect 31251 32521 31263 32524
rect 31205 32515 31263 32521
rect 32030 32512 32036 32524
rect 32088 32512 32094 32564
rect 32217 32555 32275 32561
rect 32217 32521 32229 32555
rect 32263 32552 32275 32555
rect 32306 32552 32312 32564
rect 32263 32524 32312 32552
rect 32263 32521 32275 32524
rect 32217 32515 32275 32521
rect 32306 32512 32312 32524
rect 32364 32512 32370 32564
rect 34698 32552 34704 32564
rect 32416 32524 34704 32552
rect 22097 32487 22155 32493
rect 21008 32456 21864 32484
rect 15749 32419 15807 32425
rect 15749 32385 15761 32419
rect 15795 32385 15807 32419
rect 15749 32379 15807 32385
rect 17037 32419 17095 32425
rect 17037 32385 17049 32419
rect 17083 32385 17095 32419
rect 17037 32379 17095 32385
rect 7469 32351 7527 32357
rect 7469 32348 7481 32351
rect 6604 32320 7481 32348
rect 6604 32308 6610 32320
rect 7469 32317 7481 32320
rect 7515 32317 7527 32351
rect 7469 32311 7527 32317
rect 7745 32351 7803 32357
rect 7745 32317 7757 32351
rect 7791 32348 7803 32351
rect 9858 32348 9864 32360
rect 7791 32320 9720 32348
rect 9819 32320 9864 32348
rect 7791 32317 7803 32320
rect 7745 32311 7803 32317
rect 9692 32289 9720 32320
rect 9858 32308 9864 32320
rect 9916 32308 9922 32360
rect 10321 32351 10379 32357
rect 10321 32317 10333 32351
rect 10367 32348 10379 32351
rect 10870 32348 10876 32360
rect 10367 32320 10876 32348
rect 10367 32317 10379 32320
rect 10321 32311 10379 32317
rect 9677 32283 9735 32289
rect 9677 32249 9689 32283
rect 9723 32249 9735 32283
rect 9677 32243 9735 32249
rect 1949 32215 2007 32221
rect 1949 32181 1961 32215
rect 1995 32212 2007 32215
rect 3234 32212 3240 32224
rect 1995 32184 3240 32212
rect 1995 32181 2007 32184
rect 1949 32175 2007 32181
rect 3234 32172 3240 32184
rect 3292 32172 3298 32224
rect 5718 32212 5724 32224
rect 5679 32184 5724 32212
rect 5718 32172 5724 32184
rect 5776 32172 5782 32224
rect 6825 32215 6883 32221
rect 6825 32181 6837 32215
rect 6871 32212 6883 32215
rect 8386 32212 8392 32224
rect 6871 32184 8392 32212
rect 6871 32181 6883 32184
rect 6825 32175 6883 32181
rect 8386 32172 8392 32184
rect 8444 32172 8450 32224
rect 9217 32215 9275 32221
rect 9217 32181 9229 32215
rect 9263 32212 9275 32215
rect 10336 32212 10364 32311
rect 10870 32308 10876 32320
rect 10928 32308 10934 32360
rect 12158 32348 12164 32360
rect 10980 32320 12164 32348
rect 9263 32184 10364 32212
rect 9263 32181 9275 32184
rect 9217 32175 9275 32181
rect 10410 32172 10416 32224
rect 10468 32212 10474 32224
rect 10980 32221 11008 32320
rect 12158 32308 12164 32320
rect 12216 32308 12222 32360
rect 11054 32240 11060 32292
rect 11112 32280 11118 32292
rect 15764 32280 15792 32379
rect 17218 32376 17224 32428
rect 17276 32416 17282 32428
rect 17865 32419 17923 32425
rect 17865 32416 17877 32419
rect 17276 32388 17877 32416
rect 17276 32376 17282 32388
rect 17865 32385 17877 32388
rect 17911 32385 17923 32419
rect 17865 32379 17923 32385
rect 18690 32376 18696 32428
rect 18748 32416 18754 32428
rect 18877 32419 18935 32425
rect 18877 32416 18889 32419
rect 18748 32388 18889 32416
rect 18748 32376 18754 32388
rect 18877 32385 18889 32388
rect 18923 32385 18935 32419
rect 18877 32379 18935 32385
rect 16850 32308 16856 32360
rect 16908 32348 16914 32360
rect 16945 32351 17003 32357
rect 16945 32348 16957 32351
rect 16908 32320 16957 32348
rect 16908 32308 16914 32320
rect 16945 32317 16957 32320
rect 16991 32317 17003 32351
rect 18892 32348 18920 32379
rect 19150 32376 19156 32428
rect 19208 32416 19214 32428
rect 19245 32419 19303 32425
rect 19245 32416 19257 32419
rect 19208 32388 19257 32416
rect 19208 32376 19214 32388
rect 19245 32385 19257 32388
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 19705 32419 19763 32425
rect 19705 32385 19717 32419
rect 19751 32416 19763 32419
rect 21082 32416 21088 32428
rect 19751 32388 19932 32416
rect 21043 32388 21088 32416
rect 19751 32385 19763 32388
rect 19705 32379 19763 32385
rect 19058 32348 19064 32360
rect 18892 32320 19064 32348
rect 16945 32311 17003 32317
rect 19058 32308 19064 32320
rect 19116 32308 19122 32360
rect 19334 32308 19340 32360
rect 19392 32348 19398 32360
rect 19797 32351 19855 32357
rect 19797 32348 19809 32351
rect 19392 32320 19809 32348
rect 19392 32308 19398 32320
rect 19797 32317 19809 32320
rect 19843 32317 19855 32351
rect 19797 32311 19855 32317
rect 16669 32283 16727 32289
rect 16669 32280 16681 32283
rect 11112 32252 14688 32280
rect 15764 32252 16681 32280
rect 11112 32240 11118 32252
rect 10965 32215 11023 32221
rect 10965 32212 10977 32215
rect 10468 32184 10977 32212
rect 10468 32172 10474 32184
rect 10965 32181 10977 32184
rect 11011 32181 11023 32215
rect 10965 32175 11023 32181
rect 11606 32172 11612 32224
rect 11664 32212 11670 32224
rect 13354 32212 13360 32224
rect 11664 32184 13360 32212
rect 11664 32172 11670 32184
rect 13354 32172 13360 32184
rect 13412 32172 13418 32224
rect 14660 32221 14688 32252
rect 16669 32249 16681 32252
rect 16715 32249 16727 32283
rect 16669 32243 16727 32249
rect 16758 32240 16764 32292
rect 16816 32280 16822 32292
rect 19904 32280 19932 32388
rect 21082 32376 21088 32388
rect 21140 32376 21146 32428
rect 21836 32425 21864 32456
rect 22097 32453 22109 32487
rect 22143 32453 22155 32487
rect 22097 32447 22155 32453
rect 22554 32444 22560 32496
rect 22612 32444 22618 32496
rect 24026 32444 24032 32496
rect 24084 32484 24090 32496
rect 25498 32484 25504 32496
rect 24084 32456 25504 32484
rect 24084 32444 24090 32456
rect 25498 32444 25504 32456
rect 25556 32484 25562 32496
rect 25556 32456 25636 32484
rect 25556 32444 25562 32456
rect 21821 32419 21879 32425
rect 21821 32385 21833 32419
rect 21867 32385 21879 32419
rect 24397 32419 24455 32425
rect 24397 32416 24409 32419
rect 21821 32379 21879 32385
rect 23584 32388 24409 32416
rect 23584 32360 23612 32388
rect 24397 32385 24409 32388
rect 24443 32416 24455 32419
rect 24578 32416 24584 32428
rect 24443 32388 24584 32416
rect 24443 32385 24455 32388
rect 24397 32379 24455 32385
rect 24578 32376 24584 32388
rect 24636 32376 24642 32428
rect 25608 32425 25636 32456
rect 25866 32444 25872 32496
rect 25924 32484 25930 32496
rect 26418 32484 26424 32496
rect 25924 32456 26424 32484
rect 25924 32444 25930 32456
rect 26418 32444 26424 32456
rect 26476 32484 26482 32496
rect 27985 32487 28043 32493
rect 26476 32456 27292 32484
rect 26476 32444 26482 32456
rect 25593 32419 25651 32425
rect 25593 32385 25605 32419
rect 25639 32385 25651 32419
rect 26050 32416 26056 32428
rect 26011 32388 26056 32416
rect 25593 32379 25651 32385
rect 26050 32376 26056 32388
rect 26108 32376 26114 32428
rect 26973 32419 27031 32425
rect 26973 32385 26985 32419
rect 27019 32416 27031 32419
rect 27062 32416 27068 32428
rect 27019 32388 27068 32416
rect 27019 32385 27031 32388
rect 26973 32379 27031 32385
rect 27062 32376 27068 32388
rect 27120 32376 27126 32428
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32385 27215 32419
rect 27264 32416 27292 32456
rect 27985 32453 27997 32487
rect 28031 32484 28043 32487
rect 28166 32484 28172 32496
rect 28031 32456 28172 32484
rect 28031 32453 28043 32456
rect 27985 32447 28043 32453
rect 28166 32444 28172 32456
rect 28224 32444 28230 32496
rect 28813 32487 28871 32493
rect 28813 32453 28825 32487
rect 28859 32484 28871 32487
rect 29178 32484 29184 32496
rect 28859 32456 29184 32484
rect 28859 32453 28871 32456
rect 28813 32447 28871 32453
rect 29178 32444 29184 32456
rect 29236 32444 29242 32496
rect 29730 32484 29736 32496
rect 29288 32456 29736 32484
rect 29288 32416 29316 32456
rect 29730 32444 29736 32456
rect 29788 32444 29794 32496
rect 29822 32444 29828 32496
rect 29880 32484 29886 32496
rect 30837 32487 30895 32493
rect 30837 32484 30849 32487
rect 29880 32456 30849 32484
rect 29880 32444 29886 32456
rect 30837 32453 30849 32456
rect 30883 32453 30895 32487
rect 30837 32447 30895 32453
rect 31110 32444 31116 32496
rect 31168 32484 31174 32496
rect 31168 32456 31524 32484
rect 31168 32444 31174 32456
rect 27264 32388 29316 32416
rect 29641 32419 29699 32425
rect 27157 32379 27215 32385
rect 29641 32385 29653 32419
rect 29687 32385 29699 32419
rect 29641 32379 29699 32385
rect 29917 32419 29975 32425
rect 29917 32385 29929 32419
rect 29963 32416 29975 32419
rect 30190 32416 30196 32428
rect 29963 32388 30196 32416
rect 29963 32385 29975 32388
rect 29917 32379 29975 32385
rect 23566 32348 23572 32360
rect 23479 32320 23572 32348
rect 23566 32308 23572 32320
rect 23624 32308 23630 32360
rect 24210 32348 24216 32360
rect 24171 32320 24216 32348
rect 24210 32308 24216 32320
rect 24268 32308 24274 32360
rect 24302 32308 24308 32360
rect 24360 32348 24366 32360
rect 24486 32348 24492 32360
rect 24360 32320 24405 32348
rect 24447 32320 24492 32348
rect 24360 32308 24366 32320
rect 24486 32308 24492 32320
rect 24544 32308 24550 32360
rect 25222 32308 25228 32360
rect 25280 32348 25286 32360
rect 25317 32351 25375 32357
rect 25317 32348 25329 32351
rect 25280 32320 25329 32348
rect 25280 32308 25286 32320
rect 25317 32317 25329 32320
rect 25363 32348 25375 32351
rect 25682 32348 25688 32360
rect 25363 32320 25688 32348
rect 25363 32317 25375 32320
rect 25317 32311 25375 32317
rect 25682 32308 25688 32320
rect 25740 32308 25746 32360
rect 27172 32348 27200 32379
rect 29656 32348 29684 32379
rect 30190 32376 30196 32388
rect 30248 32376 30254 32428
rect 30282 32376 30288 32428
rect 30340 32416 30346 32428
rect 31389 32419 31447 32425
rect 30340 32406 31340 32416
rect 31389 32406 31401 32419
rect 30340 32388 31401 32406
rect 30340 32376 30346 32388
rect 31312 32385 31401 32388
rect 31435 32385 31447 32419
rect 31496 32416 31524 32456
rect 31662 32444 31668 32496
rect 31720 32484 31726 32496
rect 31846 32484 31852 32496
rect 31720 32456 31852 32484
rect 31720 32444 31726 32456
rect 31846 32444 31852 32456
rect 31904 32444 31910 32496
rect 32416 32484 32444 32524
rect 34698 32512 34704 32524
rect 34756 32552 34762 32564
rect 35161 32555 35219 32561
rect 35161 32552 35173 32555
rect 34756 32524 35173 32552
rect 34756 32512 34762 32524
rect 35161 32521 35173 32524
rect 35207 32521 35219 32555
rect 37642 32552 37648 32564
rect 37603 32524 37648 32552
rect 35161 32515 35219 32521
rect 37642 32512 37648 32524
rect 37700 32512 37706 32564
rect 32232 32456 32444 32484
rect 32493 32487 32551 32493
rect 31496 32388 31984 32416
rect 31312 32379 31447 32385
rect 31312 32378 31432 32379
rect 31754 32348 31760 32360
rect 27172 32320 29592 32348
rect 29656 32320 31760 32348
rect 16816 32252 19932 32280
rect 25501 32283 25559 32289
rect 16816 32240 16822 32252
rect 25501 32249 25513 32283
rect 25547 32280 25559 32283
rect 25590 32280 25596 32292
rect 25547 32252 25596 32280
rect 25547 32249 25559 32252
rect 25501 32243 25559 32249
rect 25590 32240 25596 32252
rect 25648 32280 25654 32292
rect 27617 32283 27675 32289
rect 27617 32280 27629 32283
rect 25648 32252 27629 32280
rect 25648 32240 25654 32252
rect 27617 32249 27629 32252
rect 27663 32280 27675 32283
rect 27706 32280 27712 32292
rect 27663 32252 27712 32280
rect 27663 32249 27675 32252
rect 27617 32243 27675 32249
rect 27706 32240 27712 32252
rect 27764 32240 27770 32292
rect 28442 32280 28448 32292
rect 28355 32252 28448 32280
rect 28442 32240 28448 32252
rect 28500 32280 28506 32292
rect 29564 32280 29592 32320
rect 31754 32308 31760 32320
rect 31812 32308 31818 32360
rect 31956 32348 31984 32388
rect 32232 32348 32260 32456
rect 32493 32453 32505 32487
rect 32539 32484 32551 32487
rect 32858 32484 32864 32496
rect 32539 32456 32864 32484
rect 32539 32453 32551 32456
rect 32493 32447 32551 32453
rect 32858 32444 32864 32456
rect 32916 32444 32922 32496
rect 32398 32416 32404 32428
rect 32359 32388 32404 32416
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 32585 32419 32643 32425
rect 32585 32385 32597 32419
rect 32631 32385 32643 32419
rect 32585 32379 32643 32385
rect 32723 32419 32781 32425
rect 32723 32385 32735 32419
rect 32769 32416 32781 32419
rect 32950 32416 32956 32428
rect 32769 32388 32956 32416
rect 32769 32385 32781 32388
rect 32723 32379 32781 32385
rect 31956 32320 32260 32348
rect 32306 32308 32312 32360
rect 32364 32348 32370 32360
rect 32600 32348 32628 32379
rect 32950 32376 32956 32388
rect 33008 32376 33014 32428
rect 34790 32376 34796 32428
rect 34848 32376 34854 32428
rect 36262 32376 36268 32428
rect 36320 32416 36326 32428
rect 36541 32419 36599 32425
rect 36541 32416 36553 32419
rect 36320 32388 36553 32416
rect 36320 32376 36326 32388
rect 36541 32385 36553 32388
rect 36587 32385 36599 32419
rect 36541 32379 36599 32385
rect 37737 32419 37795 32425
rect 37737 32385 37749 32419
rect 37783 32416 37795 32419
rect 37918 32416 37924 32428
rect 37783 32388 37924 32416
rect 37783 32385 37795 32388
rect 37737 32379 37795 32385
rect 37918 32376 37924 32388
rect 37976 32376 37982 32428
rect 32364 32320 32628 32348
rect 32861 32351 32919 32357
rect 32364 32308 32370 32320
rect 32861 32317 32873 32351
rect 32907 32348 32919 32351
rect 33226 32348 33232 32360
rect 32907 32320 33232 32348
rect 32907 32317 32919 32320
rect 32861 32311 32919 32317
rect 33226 32308 33232 32320
rect 33284 32308 33290 32360
rect 33410 32348 33416 32360
rect 33371 32320 33416 32348
rect 33410 32308 33416 32320
rect 33468 32308 33474 32360
rect 33689 32351 33747 32357
rect 33689 32317 33701 32351
rect 33735 32348 33747 32351
rect 34146 32348 34152 32360
rect 33735 32320 34152 32348
rect 33735 32317 33747 32320
rect 33689 32311 33747 32317
rect 34146 32308 34152 32320
rect 34204 32308 34210 32360
rect 30742 32280 30748 32292
rect 28500 32252 28948 32280
rect 29564 32252 30748 32280
rect 28500 32240 28506 32252
rect 14645 32215 14703 32221
rect 14645 32181 14657 32215
rect 14691 32212 14703 32215
rect 18690 32212 18696 32224
rect 14691 32184 18696 32212
rect 14691 32181 14703 32184
rect 14645 32175 14703 32181
rect 18690 32172 18696 32184
rect 18748 32172 18754 32224
rect 18874 32172 18880 32224
rect 18932 32212 18938 32224
rect 19334 32212 19340 32224
rect 18932 32184 19340 32212
rect 18932 32172 18938 32184
rect 19334 32172 19340 32184
rect 19392 32172 19398 32224
rect 22094 32172 22100 32224
rect 22152 32212 22158 32224
rect 24029 32215 24087 32221
rect 24029 32212 24041 32215
rect 22152 32184 24041 32212
rect 22152 32172 22158 32184
rect 24029 32181 24041 32184
rect 24075 32181 24087 32215
rect 24029 32175 24087 32181
rect 26973 32215 27031 32221
rect 26973 32181 26985 32215
rect 27019 32212 27031 32215
rect 27338 32212 27344 32224
rect 27019 32184 27344 32212
rect 27019 32181 27031 32184
rect 26973 32175 27031 32181
rect 27338 32172 27344 32184
rect 27396 32172 27402 32224
rect 27801 32215 27859 32221
rect 27801 32181 27813 32215
rect 27847 32212 27859 32215
rect 27982 32212 27988 32224
rect 27847 32184 27988 32212
rect 27847 32181 27859 32184
rect 27801 32175 27859 32181
rect 27982 32172 27988 32184
rect 28040 32172 28046 32224
rect 28626 32212 28632 32224
rect 28587 32184 28632 32212
rect 28626 32172 28632 32184
rect 28684 32212 28690 32224
rect 28810 32212 28816 32224
rect 28684 32184 28816 32212
rect 28684 32172 28690 32184
rect 28810 32172 28816 32184
rect 28868 32172 28874 32224
rect 28920 32212 28948 32252
rect 30742 32240 30748 32252
rect 30800 32240 30806 32292
rect 31938 32280 31944 32292
rect 31496 32252 31944 32280
rect 31496 32212 31524 32252
rect 31938 32240 31944 32252
rect 31996 32240 32002 32292
rect 28920 32184 31524 32212
rect 36081 32215 36139 32221
rect 36081 32181 36093 32215
rect 36127 32212 36139 32215
rect 36262 32212 36268 32224
rect 36127 32184 36268 32212
rect 36127 32181 36139 32184
rect 36081 32175 36139 32181
rect 36262 32172 36268 32184
rect 36320 32172 36326 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 7650 31968 7656 32020
rect 7708 32008 7714 32020
rect 10597 32011 10655 32017
rect 7708 31980 9444 32008
rect 7708 31968 7714 31980
rect 7101 31943 7159 31949
rect 7101 31940 7113 31943
rect 6886 31912 7113 31940
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 3234 31872 3240 31884
rect 3195 31844 3240 31872
rect 3234 31832 3240 31844
rect 3292 31832 3298 31884
rect 6273 31875 6331 31881
rect 6273 31841 6285 31875
rect 6319 31872 6331 31875
rect 6886 31872 6914 31912
rect 7101 31909 7113 31912
rect 7147 31909 7159 31943
rect 7101 31903 7159 31909
rect 7834 31900 7840 31952
rect 7892 31940 7898 31952
rect 8389 31943 8447 31949
rect 8389 31940 8401 31943
rect 7892 31912 8401 31940
rect 7892 31900 7898 31912
rect 8389 31909 8401 31912
rect 8435 31940 8447 31943
rect 9416 31940 9444 31980
rect 10597 31977 10609 32011
rect 10643 32008 10655 32011
rect 11698 32008 11704 32020
rect 10643 31980 11704 32008
rect 10643 31977 10655 31980
rect 10597 31971 10655 31977
rect 11698 31968 11704 31980
rect 11756 31968 11762 32020
rect 11790 31968 11796 32020
rect 11848 32008 11854 32020
rect 12437 32011 12495 32017
rect 12437 32008 12449 32011
rect 11848 31980 12449 32008
rect 11848 31968 11854 31980
rect 12437 31977 12449 31980
rect 12483 31977 12495 32011
rect 12437 31971 12495 31977
rect 13170 31968 13176 32020
rect 13228 32008 13234 32020
rect 13265 32011 13323 32017
rect 13265 32008 13277 32011
rect 13228 31980 13277 32008
rect 13228 31968 13234 31980
rect 13265 31977 13277 31980
rect 13311 32008 13323 32011
rect 16758 32008 16764 32020
rect 13311 31980 16764 32008
rect 13311 31977 13323 31980
rect 13265 31971 13323 31977
rect 16758 31968 16764 31980
rect 16816 31968 16822 32020
rect 18046 31968 18052 32020
rect 18104 32008 18110 32020
rect 18509 32011 18567 32017
rect 18509 32008 18521 32011
rect 18104 31980 18521 32008
rect 18104 31968 18110 31980
rect 18509 31977 18521 31980
rect 18555 31977 18567 32011
rect 20993 32011 21051 32017
rect 20993 32008 21005 32011
rect 18509 31971 18567 31977
rect 19076 31980 21005 32008
rect 11054 31940 11060 31952
rect 8435 31912 9352 31940
rect 9416 31912 11060 31940
rect 8435 31909 8447 31912
rect 8389 31903 8447 31909
rect 7282 31872 7288 31884
rect 6319 31844 6914 31872
rect 7195 31844 7288 31872
rect 6319 31841 6331 31844
rect 6273 31835 6331 31841
rect 7282 31832 7288 31844
rect 7340 31872 7346 31884
rect 9324 31881 9352 31912
rect 11054 31900 11060 31912
rect 11112 31900 11118 31952
rect 14185 31943 14243 31949
rect 14185 31909 14197 31943
rect 14231 31940 14243 31943
rect 15286 31940 15292 31952
rect 14231 31912 15292 31940
rect 14231 31909 14243 31912
rect 14185 31903 14243 31909
rect 15286 31900 15292 31912
rect 15344 31900 15350 31952
rect 17218 31940 17224 31952
rect 17179 31912 17224 31940
rect 17218 31900 17224 31912
rect 17276 31900 17282 31952
rect 8941 31875 8999 31881
rect 8941 31872 8953 31875
rect 7340 31844 8953 31872
rect 7340 31832 7346 31844
rect 8941 31841 8953 31844
rect 8987 31841 8999 31875
rect 8941 31835 8999 31841
rect 9309 31875 9367 31881
rect 9309 31841 9321 31875
rect 9355 31841 9367 31875
rect 11333 31875 11391 31881
rect 11333 31872 11345 31875
rect 9309 31835 9367 31841
rect 10244 31844 11345 31872
rect 10244 31816 10272 31844
rect 11333 31841 11345 31844
rect 11379 31872 11391 31875
rect 11698 31872 11704 31884
rect 11379 31844 11704 31872
rect 11379 31841 11391 31844
rect 11333 31835 11391 31841
rect 11698 31832 11704 31844
rect 11756 31872 11762 31884
rect 11756 31844 12572 31872
rect 11756 31832 11762 31844
rect 6546 31764 6552 31816
rect 6604 31804 6610 31816
rect 6604 31776 6649 31804
rect 6604 31764 6610 31776
rect 7374 31764 7380 31816
rect 7432 31804 7438 31816
rect 7650 31804 7656 31816
rect 7432 31776 7477 31804
rect 7611 31776 7656 31804
rect 7432 31764 7438 31776
rect 7650 31764 7656 31776
rect 7708 31764 7714 31816
rect 7745 31807 7803 31813
rect 7745 31773 7757 31807
rect 7791 31804 7803 31807
rect 7834 31804 7840 31816
rect 7791 31776 7840 31804
rect 7791 31773 7803 31776
rect 7745 31767 7803 31773
rect 7834 31764 7840 31776
rect 7892 31764 7898 31816
rect 8205 31807 8263 31813
rect 8205 31773 8217 31807
rect 8251 31773 8263 31807
rect 8205 31767 8263 31773
rect 3050 31736 3056 31748
rect 3011 31708 3056 31736
rect 3050 31696 3056 31708
rect 3108 31696 3114 31748
rect 5718 31696 5724 31748
rect 5776 31696 5782 31748
rect 4801 31671 4859 31677
rect 4801 31637 4813 31671
rect 4847 31668 4859 31671
rect 7374 31668 7380 31680
rect 4847 31640 7380 31668
rect 4847 31637 4859 31640
rect 4801 31631 4859 31637
rect 7374 31628 7380 31640
rect 7432 31668 7438 31680
rect 8220 31668 8248 31767
rect 8294 31764 8300 31816
rect 8352 31804 8358 31816
rect 9125 31807 9183 31813
rect 9125 31804 9137 31807
rect 8352 31776 9137 31804
rect 8352 31764 8358 31776
rect 9125 31773 9137 31776
rect 9171 31804 9183 31807
rect 9858 31804 9864 31816
rect 9171 31776 9864 31804
rect 9171 31773 9183 31776
rect 9125 31767 9183 31773
rect 9858 31764 9864 31776
rect 9916 31764 9922 31816
rect 10226 31804 10232 31816
rect 10187 31776 10232 31804
rect 10226 31764 10232 31776
rect 10284 31764 10290 31816
rect 11054 31804 11060 31816
rect 10967 31776 11060 31804
rect 11054 31764 11060 31776
rect 11112 31806 11118 31816
rect 11112 31804 11192 31806
rect 11112 31778 12112 31804
rect 11112 31764 11118 31778
rect 11164 31776 12112 31778
rect 10410 31736 10416 31748
rect 10371 31708 10416 31736
rect 10410 31696 10416 31708
rect 10468 31696 10474 31748
rect 12084 31736 12112 31776
rect 12158 31764 12164 31816
rect 12216 31804 12222 31816
rect 12544 31813 12572 31844
rect 13998 31832 14004 31884
rect 14056 31872 14062 31884
rect 15565 31875 15623 31881
rect 14056 31844 15424 31872
rect 14056 31832 14062 31844
rect 12345 31807 12403 31813
rect 12345 31804 12357 31807
rect 12216 31776 12357 31804
rect 12216 31764 12222 31776
rect 12345 31773 12357 31776
rect 12391 31773 12403 31807
rect 12345 31767 12403 31773
rect 12529 31807 12587 31813
rect 12529 31773 12541 31807
rect 12575 31773 12587 31807
rect 12529 31767 12587 31773
rect 13449 31807 13507 31813
rect 13449 31773 13461 31807
rect 13495 31804 13507 31807
rect 13538 31804 13544 31816
rect 13495 31776 13544 31804
rect 13495 31773 13507 31776
rect 13449 31767 13507 31773
rect 13538 31764 13544 31776
rect 13596 31764 13602 31816
rect 14108 31813 14136 31844
rect 14093 31807 14151 31813
rect 14093 31773 14105 31807
rect 14139 31804 14151 31807
rect 14277 31807 14335 31813
rect 14139 31776 14173 31804
rect 14139 31773 14151 31776
rect 14093 31767 14151 31773
rect 14277 31773 14289 31807
rect 14323 31804 14335 31807
rect 15010 31804 15016 31816
rect 14323 31776 15016 31804
rect 14323 31773 14335 31776
rect 14277 31767 14335 31773
rect 15010 31764 15016 31776
rect 15068 31764 15074 31816
rect 15194 31764 15200 31816
rect 15252 31804 15258 31816
rect 15289 31807 15347 31813
rect 15289 31804 15301 31807
rect 15252 31776 15301 31804
rect 15252 31764 15258 31776
rect 15289 31773 15301 31776
rect 15335 31773 15347 31807
rect 15396 31804 15424 31844
rect 15565 31841 15577 31875
rect 15611 31872 15623 31875
rect 16850 31872 16856 31884
rect 15611 31844 16856 31872
rect 15611 31841 15623 31844
rect 15565 31835 15623 31841
rect 16850 31832 16856 31844
rect 16908 31832 16914 31884
rect 17773 31875 17831 31881
rect 17773 31841 17785 31875
rect 17819 31872 17831 31875
rect 18966 31872 18972 31884
rect 17819 31844 18972 31872
rect 17819 31841 17831 31844
rect 17773 31835 17831 31841
rect 18966 31832 18972 31844
rect 19024 31832 19030 31884
rect 15654 31804 15660 31816
rect 15396 31776 15660 31804
rect 15289 31767 15347 31773
rect 15654 31764 15660 31776
rect 15712 31764 15718 31816
rect 16298 31804 16304 31816
rect 16259 31776 16304 31804
rect 16298 31764 16304 31776
rect 16356 31764 16362 31816
rect 16482 31764 16488 31816
rect 16540 31804 16546 31816
rect 17037 31807 17095 31813
rect 17037 31804 17049 31807
rect 16540 31776 17049 31804
rect 16540 31764 16546 31776
rect 17037 31773 17049 31776
rect 17083 31773 17095 31807
rect 17678 31804 17684 31816
rect 17639 31776 17684 31804
rect 17037 31767 17095 31773
rect 17678 31764 17684 31776
rect 17736 31764 17742 31816
rect 17862 31804 17868 31816
rect 17823 31776 17868 31804
rect 17862 31764 17868 31776
rect 17920 31764 17926 31816
rect 13262 31736 13268 31748
rect 12084 31708 13268 31736
rect 13262 31696 13268 31708
rect 13320 31696 13326 31748
rect 18506 31745 18512 31748
rect 18493 31739 18512 31745
rect 18493 31705 18505 31739
rect 18493 31699 18512 31705
rect 18506 31696 18512 31699
rect 18564 31696 18570 31748
rect 18693 31739 18751 31745
rect 18693 31705 18705 31739
rect 18739 31736 18751 31739
rect 18782 31736 18788 31748
rect 18739 31708 18788 31736
rect 18739 31705 18751 31708
rect 18693 31699 18751 31705
rect 18782 31696 18788 31708
rect 18840 31736 18846 31748
rect 19076 31736 19104 31980
rect 20993 31977 21005 31980
rect 21039 31977 21051 32011
rect 20993 31971 21051 31977
rect 21082 31968 21088 32020
rect 21140 32008 21146 32020
rect 22557 32011 22615 32017
rect 22557 32008 22569 32011
rect 21140 31980 22569 32008
rect 21140 31968 21146 31980
rect 22557 31977 22569 31980
rect 22603 31977 22615 32011
rect 24118 32008 24124 32020
rect 22557 31971 22615 31977
rect 22848 31980 24124 32008
rect 22848 31940 22876 31980
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 24394 31968 24400 32020
rect 24452 32008 24458 32020
rect 29086 32008 29092 32020
rect 24452 31980 29092 32008
rect 24452 31968 24458 31980
rect 29086 31968 29092 31980
rect 29144 32008 29150 32020
rect 30282 32008 30288 32020
rect 29144 31980 30288 32008
rect 29144 31968 29150 31980
rect 30282 31968 30288 31980
rect 30340 31968 30346 32020
rect 31389 32011 31447 32017
rect 31389 31977 31401 32011
rect 31435 31977 31447 32011
rect 31389 31971 31447 31977
rect 21928 31912 22876 31940
rect 24949 31943 25007 31949
rect 19242 31872 19248 31884
rect 19203 31844 19248 31872
rect 19242 31832 19248 31844
rect 19300 31832 19306 31884
rect 21928 31816 21956 31912
rect 24949 31909 24961 31943
rect 24995 31940 25007 31943
rect 28166 31940 28172 31952
rect 24995 31912 28172 31940
rect 24995 31909 25007 31912
rect 24949 31903 25007 31909
rect 28166 31900 28172 31912
rect 28224 31900 28230 31952
rect 29178 31940 29184 31952
rect 29012 31912 29184 31940
rect 22005 31875 22063 31881
rect 22005 31841 22017 31875
rect 22051 31872 22063 31875
rect 22830 31872 22836 31884
rect 22051 31844 22836 31872
rect 22051 31841 22063 31844
rect 22005 31835 22063 31841
rect 22830 31832 22836 31844
rect 22888 31872 22894 31884
rect 23017 31875 23075 31881
rect 23017 31872 23029 31875
rect 22888 31844 23029 31872
rect 22888 31832 22894 31844
rect 23017 31841 23029 31844
rect 23063 31841 23075 31875
rect 23017 31835 23075 31841
rect 23201 31875 23259 31881
rect 23201 31841 23213 31875
rect 23247 31872 23259 31875
rect 23566 31872 23572 31884
rect 23247 31844 23572 31872
rect 23247 31841 23259 31844
rect 23201 31835 23259 31841
rect 23566 31832 23572 31844
rect 23624 31832 23630 31884
rect 27522 31872 27528 31884
rect 23676 31844 26372 31872
rect 20622 31764 20628 31816
rect 20680 31764 20686 31816
rect 21910 31804 21916 31816
rect 21871 31776 21916 31804
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 22094 31764 22100 31816
rect 22152 31804 22158 31816
rect 22152 31776 22197 31804
rect 22152 31764 22158 31776
rect 23382 31764 23388 31816
rect 23440 31804 23446 31816
rect 23676 31804 23704 31844
rect 23440 31776 23704 31804
rect 23440 31764 23446 31776
rect 24302 31764 24308 31816
rect 24360 31804 24366 31816
rect 24673 31807 24731 31813
rect 24673 31804 24685 31807
rect 24360 31776 24685 31804
rect 24360 31764 24366 31776
rect 24673 31773 24685 31776
rect 24719 31773 24731 31807
rect 25406 31804 25412 31816
rect 25367 31776 25412 31804
rect 24673 31767 24731 31773
rect 25406 31764 25412 31776
rect 25464 31764 25470 31816
rect 26050 31764 26056 31816
rect 26108 31804 26114 31816
rect 26145 31807 26203 31813
rect 26145 31804 26157 31807
rect 26108 31776 26157 31804
rect 26108 31764 26114 31776
rect 26145 31773 26157 31776
rect 26191 31773 26203 31807
rect 26145 31767 26203 31773
rect 18840 31708 19104 31736
rect 18840 31696 18846 31708
rect 19426 31696 19432 31748
rect 19484 31736 19490 31748
rect 19521 31739 19579 31745
rect 19521 31736 19533 31739
rect 19484 31708 19533 31736
rect 19484 31696 19490 31708
rect 19521 31705 19533 31708
rect 19567 31705 19579 31739
rect 22922 31736 22928 31748
rect 22883 31708 22928 31736
rect 19521 31699 19579 31705
rect 22922 31696 22928 31708
rect 22980 31696 22986 31748
rect 24394 31736 24400 31748
rect 24355 31708 24400 31736
rect 24394 31696 24400 31708
rect 24452 31696 24458 31748
rect 24578 31736 24584 31748
rect 24539 31708 24584 31736
rect 24578 31696 24584 31708
rect 24636 31696 24642 31748
rect 24765 31739 24823 31745
rect 24765 31705 24777 31739
rect 24811 31736 24823 31739
rect 25038 31736 25044 31748
rect 24811 31708 25044 31736
rect 24811 31705 24823 31708
rect 24765 31699 24823 31705
rect 25038 31696 25044 31708
rect 25096 31696 25102 31748
rect 7432 31640 8248 31668
rect 7432 31628 7438 31640
rect 18138 31628 18144 31680
rect 18196 31668 18202 31680
rect 18325 31671 18383 31677
rect 18325 31668 18337 31671
rect 18196 31640 18337 31668
rect 18196 31628 18202 31640
rect 18325 31637 18337 31640
rect 18371 31637 18383 31671
rect 18325 31631 18383 31637
rect 25593 31671 25651 31677
rect 25593 31637 25605 31671
rect 25639 31668 25651 31671
rect 25866 31668 25872 31680
rect 25639 31640 25872 31668
rect 25639 31637 25651 31640
rect 25593 31631 25651 31637
rect 25866 31628 25872 31640
rect 25924 31628 25930 31680
rect 26344 31677 26372 31844
rect 27356 31844 27528 31872
rect 27356 31813 27384 31844
rect 27522 31832 27528 31844
rect 27580 31832 27586 31884
rect 27982 31832 27988 31884
rect 28040 31872 28046 31884
rect 29012 31881 29040 31912
rect 29178 31900 29184 31912
rect 29236 31940 29242 31952
rect 31404 31940 31432 31971
rect 31570 31968 31576 32020
rect 31628 32008 31634 32020
rect 34606 32008 34612 32020
rect 31628 31980 34612 32008
rect 31628 31968 31634 31980
rect 34606 31968 34612 31980
rect 34664 31968 34670 32020
rect 32122 31940 32128 31952
rect 29236 31912 31432 31940
rect 31864 31912 32128 31940
rect 29236 31900 29242 31912
rect 28721 31875 28779 31881
rect 28721 31872 28733 31875
rect 28040 31844 28733 31872
rect 28040 31832 28046 31844
rect 28721 31841 28733 31844
rect 28767 31841 28779 31875
rect 28721 31835 28779 31841
rect 28997 31875 29055 31881
rect 28997 31841 29009 31875
rect 29043 31841 29055 31875
rect 29822 31872 29828 31884
rect 28997 31835 29055 31841
rect 29656 31844 29828 31872
rect 27341 31807 27399 31813
rect 27341 31773 27353 31807
rect 27387 31773 27399 31807
rect 27341 31767 27399 31773
rect 27614 31764 27620 31816
rect 27672 31804 27678 31816
rect 27709 31807 27767 31813
rect 27709 31804 27721 31807
rect 27672 31776 27721 31804
rect 27672 31764 27678 31776
rect 27709 31773 27721 31776
rect 27755 31773 27767 31807
rect 28736 31804 28764 31835
rect 29656 31804 29684 31844
rect 29822 31832 29828 31844
rect 29880 31872 29886 31884
rect 30282 31872 30288 31884
rect 29880 31844 30288 31872
rect 29880 31832 29886 31844
rect 30282 31832 30288 31844
rect 30340 31832 30346 31884
rect 30469 31875 30527 31881
rect 30469 31841 30481 31875
rect 30515 31872 30527 31875
rect 30834 31872 30840 31884
rect 30515 31844 30840 31872
rect 30515 31841 30527 31844
rect 30469 31835 30527 31841
rect 30834 31832 30840 31844
rect 30892 31832 30898 31884
rect 31864 31872 31892 31912
rect 32122 31900 32128 31912
rect 32180 31900 32186 31952
rect 32217 31943 32275 31949
rect 32217 31909 32229 31943
rect 32263 31940 32275 31943
rect 33686 31940 33692 31952
rect 32263 31912 33692 31940
rect 32263 31909 32275 31912
rect 32217 31903 32275 31909
rect 33686 31900 33692 31912
rect 33744 31900 33750 31952
rect 33796 31912 35020 31940
rect 31404 31844 31892 31872
rect 32585 31875 32643 31881
rect 28736 31776 29684 31804
rect 29733 31807 29791 31813
rect 27709 31767 27767 31773
rect 29733 31773 29745 31807
rect 29779 31804 29791 31807
rect 29914 31804 29920 31816
rect 29779 31776 29920 31804
rect 29779 31773 29791 31776
rect 29733 31767 29791 31773
rect 29914 31764 29920 31776
rect 29972 31764 29978 31816
rect 30561 31807 30619 31813
rect 30561 31773 30573 31807
rect 30607 31804 30619 31807
rect 31021 31807 31079 31813
rect 30607 31776 30972 31804
rect 30607 31773 30619 31776
rect 30561 31767 30619 31773
rect 27525 31739 27583 31745
rect 27525 31736 27537 31739
rect 26804 31708 27537 31736
rect 26804 31680 26832 31708
rect 27525 31705 27537 31708
rect 27571 31736 27583 31739
rect 27571 31708 27752 31736
rect 27571 31705 27583 31708
rect 27525 31699 27583 31705
rect 26329 31671 26387 31677
rect 26329 31637 26341 31671
rect 26375 31637 26387 31671
rect 26329 31631 26387 31637
rect 26786 31628 26792 31680
rect 26844 31628 26850 31680
rect 27724 31668 27752 31708
rect 27798 31696 27804 31748
rect 27856 31736 27862 31748
rect 30466 31736 30472 31748
rect 27856 31708 30472 31736
rect 27856 31696 27862 31708
rect 30466 31696 30472 31708
rect 30524 31696 30530 31748
rect 30944 31736 30972 31776
rect 31021 31773 31033 31807
rect 31067 31804 31079 31807
rect 31110 31804 31116 31816
rect 31067 31776 31116 31804
rect 31067 31773 31079 31776
rect 31021 31767 31079 31773
rect 31110 31764 31116 31776
rect 31168 31764 31174 31816
rect 31404 31813 31432 31844
rect 32585 31841 32597 31875
rect 32631 31872 32643 31875
rect 32950 31872 32956 31884
rect 32631 31844 32956 31872
rect 32631 31841 32643 31844
rect 32585 31835 32643 31841
rect 32950 31832 32956 31844
rect 33008 31832 33014 31884
rect 33226 31832 33232 31884
rect 33284 31872 33290 31884
rect 33505 31875 33563 31881
rect 33505 31872 33517 31875
rect 33284 31844 33517 31872
rect 33284 31832 33290 31844
rect 33505 31841 33517 31844
rect 33551 31841 33563 31875
rect 33796 31872 33824 31912
rect 34054 31872 34060 31884
rect 33505 31835 33563 31841
rect 33658 31844 33824 31872
rect 33980 31844 34060 31872
rect 31389 31807 31447 31813
rect 31389 31773 31401 31807
rect 31435 31773 31447 31807
rect 31662 31804 31668 31816
rect 31623 31776 31668 31804
rect 31389 31767 31447 31773
rect 31662 31764 31668 31776
rect 31720 31764 31726 31816
rect 31938 31764 31944 31816
rect 31996 31804 32002 31816
rect 32401 31807 32459 31813
rect 32401 31804 32413 31807
rect 31996 31776 32413 31804
rect 31996 31764 32002 31776
rect 32401 31773 32413 31776
rect 32447 31773 32459 31807
rect 32401 31767 32459 31773
rect 32490 31764 32496 31816
rect 32548 31804 32554 31816
rect 33658 31813 33686 31844
rect 33980 31813 34008 31844
rect 34054 31832 34060 31844
rect 34112 31832 34118 31884
rect 34146 31832 34152 31884
rect 34204 31872 34210 31884
rect 34698 31872 34704 31884
rect 34204 31844 34249 31872
rect 34659 31844 34704 31872
rect 34204 31832 34210 31844
rect 34698 31832 34704 31844
rect 34756 31832 34762 31884
rect 34992 31881 35020 31912
rect 34977 31875 35035 31881
rect 34977 31841 34989 31875
rect 35023 31841 35035 31875
rect 36262 31872 36268 31884
rect 36223 31844 36268 31872
rect 34977 31835 35035 31841
rect 36262 31832 36268 31844
rect 36320 31832 36326 31884
rect 33643 31807 33701 31813
rect 33643 31804 33655 31807
rect 32548 31776 33655 31804
rect 32548 31764 32554 31776
rect 33643 31773 33655 31776
rect 33689 31773 33701 31807
rect 33643 31767 33701 31773
rect 33965 31807 34023 31813
rect 33965 31773 33977 31807
rect 34011 31773 34023 31807
rect 38102 31804 38108 31816
rect 38063 31776 38108 31804
rect 33965 31767 34023 31773
rect 38102 31764 38108 31776
rect 38160 31764 38166 31816
rect 31570 31736 31576 31748
rect 30944 31708 31576 31736
rect 31570 31696 31576 31708
rect 31628 31696 31634 31748
rect 33778 31736 33784 31748
rect 33739 31708 33784 31736
rect 33778 31696 33784 31708
rect 33836 31696 33842 31748
rect 33870 31696 33876 31748
rect 33928 31736 33934 31748
rect 36446 31736 36452 31748
rect 33928 31708 33973 31736
rect 36407 31708 36452 31736
rect 33928 31696 33934 31708
rect 36446 31696 36452 31708
rect 36504 31696 36510 31748
rect 28350 31668 28356 31680
rect 27724 31640 28356 31668
rect 28350 31628 28356 31640
rect 28408 31628 28414 31680
rect 29825 31671 29883 31677
rect 29825 31637 29837 31671
rect 29871 31668 29883 31671
rect 29914 31668 29920 31680
rect 29871 31640 29920 31668
rect 29871 31637 29883 31640
rect 29825 31631 29883 31637
rect 29914 31628 29920 31640
rect 29972 31628 29978 31680
rect 30006 31628 30012 31680
rect 30064 31668 30070 31680
rect 31205 31671 31263 31677
rect 31205 31668 31217 31671
rect 30064 31640 31217 31668
rect 30064 31628 30070 31640
rect 31205 31637 31217 31640
rect 31251 31637 31263 31671
rect 31205 31631 31263 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 2133 31467 2191 31473
rect 2133 31433 2145 31467
rect 2179 31464 2191 31467
rect 3050 31464 3056 31476
rect 2179 31436 3056 31464
rect 2179 31433 2191 31436
rect 2133 31427 2191 31433
rect 3050 31424 3056 31436
rect 3108 31424 3114 31476
rect 5721 31467 5779 31473
rect 5721 31433 5733 31467
rect 5767 31464 5779 31467
rect 6822 31464 6828 31476
rect 5767 31436 6828 31464
rect 5767 31433 5779 31436
rect 5721 31427 5779 31433
rect 6822 31424 6828 31436
rect 6880 31424 6886 31476
rect 7742 31424 7748 31476
rect 7800 31464 7806 31476
rect 7800 31436 7880 31464
rect 7800 31424 7806 31436
rect 7282 31396 7288 31408
rect 5828 31368 7288 31396
rect 2225 31331 2283 31337
rect 2225 31297 2237 31331
rect 2271 31328 2283 31331
rect 2314 31328 2320 31340
rect 2271 31300 2320 31328
rect 2271 31297 2283 31300
rect 2225 31291 2283 31297
rect 2314 31288 2320 31300
rect 2372 31288 2378 31340
rect 5828 31337 5856 31368
rect 7282 31356 7288 31368
rect 7340 31356 7346 31408
rect 7653 31399 7711 31405
rect 7653 31396 7665 31399
rect 7392 31368 7665 31396
rect 5169 31331 5227 31337
rect 5169 31297 5181 31331
rect 5215 31297 5227 31331
rect 5169 31291 5227 31297
rect 5629 31331 5687 31337
rect 5629 31297 5641 31331
rect 5675 31297 5687 31331
rect 5629 31291 5687 31297
rect 5813 31331 5871 31337
rect 5813 31297 5825 31331
rect 5859 31297 5871 31331
rect 5813 31291 5871 31297
rect 5184 31136 5212 31291
rect 5644 31192 5672 31291
rect 5902 31288 5908 31340
rect 5960 31328 5966 31340
rect 6641 31331 6699 31337
rect 6641 31328 6653 31331
rect 5960 31300 6653 31328
rect 5960 31288 5966 31300
rect 6641 31297 6653 31300
rect 6687 31297 6699 31331
rect 7392 31328 7420 31368
rect 7653 31365 7665 31368
rect 7699 31365 7711 31399
rect 7653 31359 7711 31365
rect 7742 31328 7748 31340
rect 6641 31291 6699 31297
rect 6840 31300 7420 31328
rect 7703 31300 7748 31328
rect 6840 31201 6868 31300
rect 7300 31272 7328 31300
rect 7742 31288 7748 31300
rect 7800 31288 7806 31340
rect 7852 31337 7880 31436
rect 9858 31424 9864 31476
rect 9916 31464 9922 31476
rect 10229 31467 10287 31473
rect 10229 31464 10241 31467
rect 9916 31436 10241 31464
rect 9916 31424 9922 31436
rect 10229 31433 10241 31436
rect 10275 31433 10287 31467
rect 10229 31427 10287 31433
rect 10397 31467 10455 31473
rect 10397 31433 10409 31467
rect 10443 31464 10455 31467
rect 11054 31464 11060 31476
rect 10443 31436 11060 31464
rect 10443 31433 10455 31436
rect 10397 31427 10455 31433
rect 11054 31424 11060 31436
rect 11112 31424 11118 31476
rect 16022 31424 16028 31476
rect 16080 31464 16086 31476
rect 16390 31464 16396 31476
rect 16080 31436 16396 31464
rect 16080 31424 16086 31436
rect 16390 31424 16396 31436
rect 16448 31424 16454 31476
rect 17678 31464 17684 31476
rect 17639 31436 17684 31464
rect 17678 31424 17684 31436
rect 17736 31424 17742 31476
rect 18138 31424 18144 31476
rect 18196 31464 18202 31476
rect 19058 31464 19064 31476
rect 18196 31436 19064 31464
rect 18196 31424 18202 31436
rect 19058 31424 19064 31436
rect 19116 31424 19122 31476
rect 19245 31467 19303 31473
rect 19245 31433 19257 31467
rect 19291 31464 19303 31467
rect 19426 31464 19432 31476
rect 19291 31436 19432 31464
rect 19291 31433 19303 31436
rect 19245 31427 19303 31433
rect 19426 31424 19432 31436
rect 19484 31424 19490 31476
rect 20622 31464 20628 31476
rect 20583 31436 20628 31464
rect 20622 31424 20628 31436
rect 20680 31424 20686 31476
rect 22281 31467 22339 31473
rect 22281 31433 22293 31467
rect 22327 31464 22339 31467
rect 22554 31464 22560 31476
rect 22327 31436 22560 31464
rect 22327 31433 22339 31436
rect 22281 31427 22339 31433
rect 22554 31424 22560 31436
rect 22612 31424 22618 31476
rect 22830 31424 22836 31476
rect 22888 31464 22894 31476
rect 23293 31467 23351 31473
rect 23293 31464 23305 31467
rect 22888 31436 23305 31464
rect 22888 31424 22894 31436
rect 23293 31433 23305 31436
rect 23339 31433 23351 31467
rect 24210 31464 24216 31476
rect 24171 31436 24216 31464
rect 23293 31427 23351 31433
rect 24210 31424 24216 31436
rect 24268 31424 24274 31476
rect 24302 31424 24308 31476
rect 24360 31464 24366 31476
rect 24397 31467 24455 31473
rect 24397 31464 24409 31467
rect 24360 31436 24409 31464
rect 24360 31424 24366 31436
rect 24397 31433 24409 31436
rect 24443 31433 24455 31467
rect 24397 31427 24455 31433
rect 25225 31467 25283 31473
rect 25225 31433 25237 31467
rect 25271 31464 25283 31467
rect 25314 31464 25320 31476
rect 25271 31436 25320 31464
rect 25271 31433 25283 31436
rect 25225 31427 25283 31433
rect 25314 31424 25320 31436
rect 25372 31464 25378 31476
rect 27798 31464 27804 31476
rect 25372 31436 27804 31464
rect 25372 31424 25378 31436
rect 27798 31424 27804 31436
rect 27856 31424 27862 31476
rect 28966 31436 30328 31464
rect 9401 31399 9459 31405
rect 9401 31365 9413 31399
rect 9447 31365 9459 31399
rect 9401 31359 9459 31365
rect 7837 31331 7895 31337
rect 7837 31297 7849 31331
rect 7883 31328 7895 31331
rect 7926 31328 7932 31340
rect 7883 31300 7932 31328
rect 7883 31297 7895 31300
rect 7837 31291 7895 31297
rect 7926 31288 7932 31300
rect 7984 31328 7990 31340
rect 8202 31328 8208 31340
rect 7984 31300 8208 31328
rect 7984 31288 7990 31300
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 8941 31331 8999 31337
rect 8941 31297 8953 31331
rect 8987 31297 8999 31331
rect 9416 31328 9444 31359
rect 9490 31356 9496 31408
rect 9548 31396 9554 31408
rect 9601 31399 9659 31405
rect 9601 31396 9613 31399
rect 9548 31368 9613 31396
rect 9548 31356 9554 31368
rect 9601 31365 9613 31368
rect 9647 31365 9659 31399
rect 9601 31359 9659 31365
rect 10597 31399 10655 31405
rect 10597 31365 10609 31399
rect 10643 31396 10655 31399
rect 10870 31396 10876 31408
rect 10643 31368 10876 31396
rect 10643 31365 10655 31368
rect 10597 31359 10655 31365
rect 10042 31328 10048 31340
rect 9416 31300 10048 31328
rect 8941 31291 8999 31297
rect 7282 31220 7288 31272
rect 7340 31220 7346 31272
rect 6825 31195 6883 31201
rect 6825 31192 6837 31195
rect 5644 31164 6837 31192
rect 6825 31161 6837 31164
rect 6871 31161 6883 31195
rect 7466 31192 7472 31204
rect 7427 31164 7472 31192
rect 6825 31155 6883 31161
rect 7466 31152 7472 31164
rect 7524 31152 7530 31204
rect 8757 31195 8815 31201
rect 8757 31192 8769 31195
rect 7576 31164 8769 31192
rect 5074 31124 5080 31136
rect 5035 31096 5080 31124
rect 5074 31084 5080 31096
rect 5132 31084 5138 31136
rect 5166 31084 5172 31136
rect 5224 31124 5230 31136
rect 6730 31124 6736 31136
rect 5224 31096 6736 31124
rect 5224 31084 5230 31096
rect 6730 31084 6736 31096
rect 6788 31124 6794 31136
rect 7576 31124 7604 31164
rect 8757 31161 8769 31164
rect 8803 31161 8815 31195
rect 8956 31192 8984 31291
rect 10042 31288 10048 31300
rect 10100 31288 10106 31340
rect 10226 31288 10232 31340
rect 10284 31328 10290 31340
rect 10612 31328 10640 31359
rect 10870 31356 10876 31368
rect 10928 31356 10934 31408
rect 11514 31396 11520 31408
rect 11475 31368 11520 31396
rect 11514 31356 11520 31368
rect 11572 31356 11578 31408
rect 11717 31399 11775 31405
rect 11717 31396 11729 31399
rect 11624 31368 11729 31396
rect 10284 31300 10640 31328
rect 10284 31288 10290 31300
rect 11624 31272 11652 31368
rect 11717 31365 11729 31368
rect 11763 31365 11775 31399
rect 14274 31396 14280 31408
rect 13846 31368 14280 31396
rect 11717 31359 11775 31365
rect 14274 31356 14280 31368
rect 14332 31356 14338 31408
rect 14737 31399 14795 31405
rect 14737 31365 14749 31399
rect 14783 31396 14795 31399
rect 16482 31396 16488 31408
rect 14783 31368 16488 31396
rect 14783 31365 14795 31368
rect 14737 31359 14795 31365
rect 16482 31356 16488 31368
rect 16540 31356 16546 31408
rect 18414 31356 18420 31408
rect 18472 31396 18478 31408
rect 19797 31399 19855 31405
rect 19797 31396 19809 31399
rect 18472 31368 19809 31396
rect 18472 31356 18478 31368
rect 19797 31365 19809 31368
rect 19843 31365 19855 31399
rect 23382 31396 23388 31408
rect 19797 31359 19855 31365
rect 22388 31368 23388 31396
rect 12342 31328 12348 31340
rect 12303 31300 12348 31328
rect 12342 31288 12348 31300
rect 12400 31288 12406 31340
rect 15010 31288 15016 31340
rect 15068 31328 15074 31340
rect 15473 31331 15531 31337
rect 15473 31328 15485 31331
rect 15068 31300 15485 31328
rect 15068 31288 15074 31300
rect 15473 31297 15485 31300
rect 15519 31297 15531 31331
rect 15473 31291 15531 31297
rect 15654 31288 15660 31340
rect 15712 31328 15718 31340
rect 16390 31328 16396 31340
rect 15712 31300 16396 31328
rect 15712 31288 15718 31300
rect 16390 31288 16396 31300
rect 16448 31288 16454 31340
rect 16574 31288 16580 31340
rect 16632 31328 16638 31340
rect 17129 31331 17187 31337
rect 17129 31328 17141 31331
rect 16632 31300 17141 31328
rect 16632 31288 16638 31300
rect 17129 31297 17141 31300
rect 17175 31328 17187 31331
rect 17402 31328 17408 31340
rect 17175 31300 17408 31328
rect 17175 31297 17187 31300
rect 17129 31291 17187 31297
rect 17402 31288 17408 31300
rect 17460 31288 17466 31340
rect 17865 31331 17923 31337
rect 17865 31297 17877 31331
rect 17911 31297 17923 31331
rect 18046 31328 18052 31340
rect 18007 31300 18052 31328
rect 17865 31291 17923 31297
rect 11606 31260 11612 31272
rect 9784 31232 11612 31260
rect 9784 31201 9812 31232
rect 11606 31220 11612 31232
rect 11664 31220 11670 31272
rect 12621 31263 12679 31269
rect 12621 31229 12633 31263
rect 12667 31260 12679 31263
rect 12710 31260 12716 31272
rect 12667 31232 12716 31260
rect 12667 31229 12679 31232
rect 12621 31223 12679 31229
rect 12710 31220 12716 31232
rect 12768 31220 12774 31272
rect 12986 31220 12992 31272
rect 13044 31260 13050 31272
rect 17880 31260 17908 31291
rect 18046 31288 18052 31300
rect 18104 31288 18110 31340
rect 18138 31288 18144 31340
rect 18196 31328 18202 31340
rect 18506 31328 18512 31340
rect 18196 31300 18512 31328
rect 18196 31288 18202 31300
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 18601 31331 18659 31337
rect 18601 31297 18613 31331
rect 18647 31328 18659 31331
rect 18782 31328 18788 31340
rect 18647 31300 18788 31328
rect 18647 31297 18659 31300
rect 18601 31291 18659 31297
rect 18414 31260 18420 31272
rect 13044 31232 16160 31260
rect 17880 31232 18420 31260
rect 13044 31220 13050 31232
rect 16132 31204 16160 31232
rect 18414 31220 18420 31232
rect 18472 31260 18478 31272
rect 18616 31260 18644 31291
rect 18782 31288 18788 31300
rect 18840 31288 18846 31340
rect 18966 31328 18972 31340
rect 18927 31300 18972 31328
rect 18966 31288 18972 31300
rect 19024 31288 19030 31340
rect 19058 31288 19064 31340
rect 19116 31328 19122 31340
rect 19889 31331 19947 31337
rect 19116 31300 19161 31328
rect 19116 31288 19122 31300
rect 19889 31297 19901 31331
rect 19935 31328 19947 31331
rect 19978 31328 19984 31340
rect 19935 31300 19984 31328
rect 19935 31297 19947 31300
rect 19889 31291 19947 31297
rect 19978 31288 19984 31300
rect 20036 31328 20042 31340
rect 20162 31328 20168 31340
rect 20036 31300 20168 31328
rect 20036 31288 20042 31300
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 20714 31328 20720 31340
rect 20675 31300 20720 31328
rect 20714 31288 20720 31300
rect 20772 31288 20778 31340
rect 22388 31337 22416 31368
rect 23382 31356 23388 31368
rect 23440 31356 23446 31408
rect 24578 31396 24584 31408
rect 24539 31368 24584 31396
rect 24578 31356 24584 31368
rect 24636 31356 24642 31408
rect 25406 31396 25412 31408
rect 24872 31368 25412 31396
rect 22373 31331 22431 31337
rect 22373 31297 22385 31331
rect 22419 31297 22431 31331
rect 22373 31291 22431 31297
rect 23201 31331 23259 31337
rect 23201 31297 23213 31331
rect 23247 31328 23259 31331
rect 24029 31331 24087 31337
rect 24029 31328 24041 31331
rect 23247 31300 24041 31328
rect 23247 31297 23259 31300
rect 23201 31291 23259 31297
rect 24029 31297 24041 31300
rect 24075 31297 24087 31331
rect 24029 31291 24087 31297
rect 24305 31331 24363 31337
rect 24305 31297 24317 31331
rect 24351 31328 24363 31331
rect 24872 31328 24900 31368
rect 25406 31356 25412 31368
rect 25464 31356 25470 31408
rect 26973 31399 27031 31405
rect 26973 31365 26985 31399
rect 27019 31396 27031 31399
rect 27062 31396 27068 31408
rect 27019 31368 27068 31396
rect 27019 31365 27031 31368
rect 26973 31359 27031 31365
rect 27062 31356 27068 31368
rect 27120 31356 27126 31408
rect 24351 31300 24900 31328
rect 24351 31297 24363 31300
rect 24305 31291 24363 31297
rect 25038 31288 25044 31340
rect 25096 31328 25102 31340
rect 26050 31328 26056 31340
rect 25096 31300 26056 31328
rect 25096 31288 25102 31300
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31328 26387 31331
rect 26510 31328 26516 31340
rect 26375 31300 26516 31328
rect 26375 31297 26387 31300
rect 26329 31291 26387 31297
rect 26510 31288 26516 31300
rect 26568 31288 26574 31340
rect 26602 31288 26608 31340
rect 26660 31328 26666 31340
rect 27157 31331 27215 31337
rect 27157 31328 27169 31331
rect 26660 31300 27169 31328
rect 26660 31288 26666 31300
rect 27157 31297 27169 31300
rect 27203 31328 27215 31331
rect 27985 31331 28043 31337
rect 27985 31328 27997 31331
rect 27203 31300 27997 31328
rect 27203 31297 27215 31300
rect 27157 31291 27215 31297
rect 27985 31297 27997 31300
rect 28031 31297 28043 31331
rect 28350 31328 28356 31340
rect 28311 31300 28356 31328
rect 27985 31291 28043 31297
rect 28350 31288 28356 31300
rect 28408 31288 28414 31340
rect 18472 31232 18644 31260
rect 18472 31220 18478 31232
rect 18690 31220 18696 31272
rect 18748 31260 18754 31272
rect 20898 31260 20904 31272
rect 18748 31232 20904 31260
rect 18748 31220 18754 31232
rect 20898 31220 20904 31232
rect 20956 31220 20962 31272
rect 23477 31263 23535 31269
rect 23477 31229 23489 31263
rect 23523 31260 23535 31263
rect 23658 31260 23664 31272
rect 23523 31232 23664 31260
rect 23523 31229 23535 31232
rect 23477 31223 23535 31229
rect 23658 31220 23664 31232
rect 23716 31260 23722 31272
rect 24394 31260 24400 31272
rect 23716 31232 24400 31260
rect 23716 31220 23722 31232
rect 24394 31220 24400 31232
rect 24452 31220 24458 31272
rect 27893 31263 27951 31269
rect 27893 31229 27905 31263
rect 27939 31260 27951 31263
rect 28718 31260 28724 31272
rect 27939 31232 28724 31260
rect 27939 31229 27951 31232
rect 27893 31223 27951 31229
rect 28718 31220 28724 31232
rect 28776 31220 28782 31272
rect 9769 31195 9827 31201
rect 8956 31164 9720 31192
rect 8757 31155 8815 31161
rect 6788 31096 7604 31124
rect 8021 31127 8079 31133
rect 6788 31084 6794 31096
rect 8021 31093 8033 31127
rect 8067 31124 8079 31127
rect 8294 31124 8300 31136
rect 8067 31096 8300 31124
rect 8067 31093 8079 31096
rect 8021 31087 8079 31093
rect 8294 31084 8300 31096
rect 8352 31084 8358 31136
rect 9582 31124 9588 31136
rect 9543 31096 9588 31124
rect 9582 31084 9588 31096
rect 9640 31084 9646 31136
rect 9692 31124 9720 31164
rect 9769 31161 9781 31195
rect 9815 31161 9827 31195
rect 9769 31155 9827 31161
rect 14366 31152 14372 31204
rect 14424 31192 14430 31204
rect 14550 31192 14556 31204
rect 14424 31164 14556 31192
rect 14424 31152 14430 31164
rect 14550 31152 14556 31164
rect 14608 31152 14614 31204
rect 16114 31152 16120 31204
rect 16172 31192 16178 31204
rect 16945 31195 17003 31201
rect 16945 31192 16957 31195
rect 16172 31164 16957 31192
rect 16172 31152 16178 31164
rect 16945 31161 16957 31164
rect 16991 31161 17003 31195
rect 16945 31155 17003 31161
rect 22002 31152 22008 31204
rect 22060 31192 22066 31204
rect 25866 31192 25872 31204
rect 22060 31164 25872 31192
rect 22060 31152 22066 31164
rect 25866 31152 25872 31164
rect 25924 31152 25930 31204
rect 26142 31192 26148 31204
rect 26103 31164 26148 31192
rect 26142 31152 26148 31164
rect 26200 31152 26206 31204
rect 28966 31192 28994 31436
rect 29914 31356 29920 31408
rect 29972 31356 29978 31408
rect 30300 31396 30328 31436
rect 30374 31424 30380 31476
rect 30432 31464 30438 31476
rect 30432 31436 31432 31464
rect 30432 31424 30438 31436
rect 30650 31396 30656 31408
rect 30300 31368 30656 31396
rect 30650 31356 30656 31368
rect 30708 31396 30714 31408
rect 30708 31368 31202 31396
rect 30708 31356 30714 31368
rect 30650 31260 30656 31272
rect 30611 31232 30656 31260
rect 30650 31220 30656 31232
rect 30708 31220 30714 31272
rect 30926 31260 30932 31272
rect 30887 31232 30932 31260
rect 30926 31220 30932 31232
rect 30984 31220 30990 31272
rect 31174 31260 31202 31368
rect 31404 31337 31432 31436
rect 31754 31424 31760 31476
rect 31812 31464 31818 31476
rect 32125 31467 32183 31473
rect 32125 31464 32137 31467
rect 31812 31436 32137 31464
rect 31812 31424 31818 31436
rect 32125 31433 32137 31436
rect 32171 31433 32183 31467
rect 32125 31427 32183 31433
rect 32858 31424 32864 31476
rect 32916 31464 32922 31476
rect 32953 31467 33011 31473
rect 32953 31464 32965 31467
rect 32916 31436 32965 31464
rect 32916 31424 32922 31436
rect 32953 31433 32965 31436
rect 32999 31433 33011 31467
rect 33870 31464 33876 31476
rect 33831 31436 33876 31464
rect 32953 31427 33011 31433
rect 33870 31424 33876 31436
rect 33928 31424 33934 31476
rect 36446 31424 36452 31476
rect 36504 31464 36510 31476
rect 36633 31467 36691 31473
rect 36633 31464 36645 31467
rect 36504 31436 36645 31464
rect 36504 31424 36510 31436
rect 36633 31433 36645 31436
rect 36679 31433 36691 31467
rect 36633 31427 36691 31433
rect 32217 31399 32275 31405
rect 32217 31365 32229 31399
rect 32263 31396 32275 31399
rect 32490 31396 32496 31408
rect 32263 31368 32496 31396
rect 32263 31365 32275 31368
rect 32217 31359 32275 31365
rect 32490 31356 32496 31368
rect 32548 31396 32554 31408
rect 32548 31368 34008 31396
rect 32548 31356 32554 31368
rect 31389 31331 31447 31337
rect 31389 31297 31401 31331
rect 31435 31297 31447 31331
rect 31389 31291 31447 31297
rect 31478 31288 31484 31340
rect 31536 31328 31542 31340
rect 31573 31331 31631 31337
rect 31573 31328 31585 31331
rect 31536 31300 31585 31328
rect 31536 31288 31542 31300
rect 31573 31297 31585 31300
rect 31619 31297 31631 31331
rect 31573 31291 31631 31297
rect 32125 31331 32183 31337
rect 32125 31297 32137 31331
rect 32171 31297 32183 31331
rect 32125 31291 32183 31297
rect 32401 31331 32459 31337
rect 32401 31297 32413 31331
rect 32447 31328 32459 31331
rect 33045 31331 33103 31337
rect 33045 31328 33057 31331
rect 32447 31300 33057 31328
rect 32447 31297 32459 31300
rect 32401 31291 32459 31297
rect 33045 31297 33057 31300
rect 33091 31328 33103 31331
rect 33686 31328 33692 31340
rect 33091 31300 33692 31328
rect 33091 31297 33103 31300
rect 33045 31291 33103 31297
rect 32140 31260 32168 31291
rect 33686 31288 33692 31300
rect 33744 31328 33750 31340
rect 33980 31337 34008 31368
rect 33781 31331 33839 31337
rect 33781 31328 33793 31331
rect 33744 31300 33793 31328
rect 33744 31288 33750 31300
rect 33781 31297 33793 31300
rect 33827 31297 33839 31331
rect 33781 31291 33839 31297
rect 33965 31331 34023 31337
rect 33965 31297 33977 31331
rect 34011 31297 34023 31331
rect 34606 31328 34612 31340
rect 34567 31300 34612 31328
rect 33965 31291 34023 31297
rect 34606 31288 34612 31300
rect 34664 31288 34670 31340
rect 36725 31331 36783 31337
rect 36725 31297 36737 31331
rect 36771 31328 36783 31331
rect 36906 31328 36912 31340
rect 36771 31300 36912 31328
rect 36771 31297 36783 31300
rect 36725 31291 36783 31297
rect 36906 31288 36912 31300
rect 36964 31288 36970 31340
rect 37645 31331 37703 31337
rect 37645 31297 37657 31331
rect 37691 31328 37703 31331
rect 37918 31328 37924 31340
rect 37691 31300 37924 31328
rect 37691 31297 37703 31300
rect 37645 31291 37703 31297
rect 37918 31288 37924 31300
rect 37976 31288 37982 31340
rect 31174 31232 32168 31260
rect 28368 31164 28994 31192
rect 10134 31124 10140 31136
rect 9692 31096 10140 31124
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 10410 31124 10416 31136
rect 10371 31096 10416 31124
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 11698 31124 11704 31136
rect 11659 31096 11704 31124
rect 11698 31084 11704 31096
rect 11756 31084 11762 31136
rect 11885 31127 11943 31133
rect 11885 31093 11897 31127
rect 11931 31124 11943 31127
rect 12158 31124 12164 31136
rect 11931 31096 12164 31124
rect 11931 31093 11943 31096
rect 11885 31087 11943 31093
rect 12158 31084 12164 31096
rect 12216 31084 12222 31136
rect 12342 31084 12348 31136
rect 12400 31124 12406 31136
rect 13354 31124 13360 31136
rect 12400 31096 13360 31124
rect 12400 31084 12406 31096
rect 13354 31084 13360 31096
rect 13412 31124 13418 31136
rect 14093 31127 14151 31133
rect 14093 31124 14105 31127
rect 13412 31096 14105 31124
rect 13412 31084 13418 31096
rect 14093 31093 14105 31096
rect 14139 31093 14151 31127
rect 14093 31087 14151 31093
rect 15289 31127 15347 31133
rect 15289 31093 15301 31127
rect 15335 31124 15347 31127
rect 15470 31124 15476 31136
rect 15335 31096 15476 31124
rect 15335 31093 15347 31096
rect 15289 31087 15347 31093
rect 15470 31084 15476 31096
rect 15528 31084 15534 31136
rect 22554 31084 22560 31136
rect 22612 31124 22618 31136
rect 22833 31127 22891 31133
rect 22833 31124 22845 31127
rect 22612 31096 22845 31124
rect 22612 31084 22618 31096
rect 22833 31093 22845 31096
rect 22879 31093 22891 31127
rect 22833 31087 22891 31093
rect 27154 31084 27160 31136
rect 27212 31124 27218 31136
rect 28368 31133 28396 31164
rect 31110 31152 31116 31204
rect 31168 31192 31174 31204
rect 32306 31192 32312 31204
rect 31168 31164 32312 31192
rect 31168 31152 31174 31164
rect 32306 31152 32312 31164
rect 32364 31152 32370 31204
rect 27341 31127 27399 31133
rect 27341 31124 27353 31127
rect 27212 31096 27353 31124
rect 27212 31084 27218 31096
rect 27341 31093 27353 31096
rect 27387 31093 27399 31127
rect 27341 31087 27399 31093
rect 28353 31127 28411 31133
rect 28353 31093 28365 31127
rect 28399 31093 28411 31127
rect 28534 31124 28540 31136
rect 28495 31096 28540 31124
rect 28353 31087 28411 31093
rect 28534 31084 28540 31096
rect 28592 31084 28598 31136
rect 29178 31124 29184 31136
rect 29139 31096 29184 31124
rect 29178 31084 29184 31096
rect 29236 31084 29242 31136
rect 29914 31084 29920 31136
rect 29972 31124 29978 31136
rect 31573 31127 31631 31133
rect 31573 31124 31585 31127
rect 29972 31096 31585 31124
rect 29972 31084 29978 31096
rect 31573 31093 31585 31096
rect 31619 31093 31631 31127
rect 31573 31087 31631 31093
rect 33042 31084 33048 31136
rect 33100 31124 33106 31136
rect 34517 31127 34575 31133
rect 34517 31124 34529 31127
rect 33100 31096 34529 31124
rect 33100 31084 33106 31096
rect 34517 31093 34529 31096
rect 34563 31093 34575 31127
rect 35434 31124 35440 31136
rect 35395 31096 35440 31124
rect 34517 31087 34575 31093
rect 35434 31084 35440 31096
rect 35492 31084 35498 31136
rect 36078 31124 36084 31136
rect 36039 31096 36084 31124
rect 36078 31084 36084 31096
rect 36136 31084 36142 31136
rect 36446 31084 36452 31136
rect 36504 31124 36510 31136
rect 37553 31127 37611 31133
rect 37553 31124 37565 31127
rect 36504 31096 37565 31124
rect 36504 31084 36510 31096
rect 37553 31093 37565 31096
rect 37599 31093 37611 31127
rect 37553 31087 37611 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 7742 30880 7748 30932
rect 7800 30920 7806 30932
rect 8205 30923 8263 30929
rect 8205 30920 8217 30923
rect 7800 30892 8217 30920
rect 7800 30880 7806 30892
rect 8205 30889 8217 30892
rect 8251 30889 8263 30923
rect 9490 30920 9496 30932
rect 9451 30892 9496 30920
rect 8205 30883 8263 30889
rect 9490 30880 9496 30892
rect 9548 30880 9554 30932
rect 9677 30923 9735 30929
rect 9677 30889 9689 30923
rect 9723 30920 9735 30923
rect 10226 30920 10232 30932
rect 9723 30892 10232 30920
rect 9723 30889 9735 30892
rect 9677 30883 9735 30889
rect 10226 30880 10232 30892
rect 10284 30880 10290 30932
rect 10594 30920 10600 30932
rect 10555 30892 10600 30920
rect 10594 30880 10600 30892
rect 10652 30880 10658 30932
rect 11057 30923 11115 30929
rect 11057 30889 11069 30923
rect 11103 30920 11115 30923
rect 17954 30920 17960 30932
rect 11103 30892 17960 30920
rect 11103 30889 11115 30892
rect 11057 30883 11115 30889
rect 17954 30880 17960 30892
rect 18012 30880 18018 30932
rect 19978 30880 19984 30932
rect 20036 30920 20042 30932
rect 23474 30920 23480 30932
rect 20036 30892 23480 30920
rect 20036 30880 20042 30892
rect 23474 30880 23480 30892
rect 23532 30880 23538 30932
rect 23658 30920 23664 30932
rect 23619 30892 23664 30920
rect 23658 30880 23664 30892
rect 23716 30880 23722 30932
rect 25866 30880 25872 30932
rect 25924 30920 25930 30932
rect 29549 30923 29607 30929
rect 25924 30892 27108 30920
rect 25924 30880 25930 30892
rect 7561 30855 7619 30861
rect 7561 30821 7573 30855
rect 7607 30852 7619 30855
rect 9582 30852 9588 30864
rect 7607 30824 9588 30852
rect 7607 30821 7619 30824
rect 7561 30815 7619 30821
rect 9582 30812 9588 30824
rect 9640 30812 9646 30864
rect 11698 30852 11704 30864
rect 11532 30824 11704 30852
rect 6089 30787 6147 30793
rect 6089 30753 6101 30787
rect 6135 30784 6147 30787
rect 6546 30784 6552 30796
rect 6135 30756 6552 30784
rect 6135 30753 6147 30756
rect 6089 30747 6147 30753
rect 6546 30744 6552 30756
rect 6604 30744 6610 30796
rect 7006 30744 7012 30796
rect 7064 30784 7070 30796
rect 7834 30784 7840 30796
rect 7064 30756 7840 30784
rect 7064 30744 7070 30756
rect 7834 30744 7840 30756
rect 7892 30744 7898 30796
rect 10778 30784 10784 30796
rect 10739 30756 10784 30784
rect 10778 30744 10784 30756
rect 10836 30744 10842 30796
rect 11532 30793 11560 30824
rect 11698 30812 11704 30824
rect 11756 30812 11762 30864
rect 14090 30852 14096 30864
rect 12544 30824 14096 30852
rect 11517 30787 11575 30793
rect 11517 30753 11529 30787
rect 11563 30753 11575 30787
rect 11517 30747 11575 30753
rect 7193 30719 7251 30725
rect 7193 30685 7205 30719
rect 7239 30716 7251 30719
rect 7466 30716 7472 30728
rect 7239 30688 7472 30716
rect 7239 30685 7251 30688
rect 7193 30679 7251 30685
rect 7466 30676 7472 30688
rect 7524 30676 7530 30728
rect 8018 30716 8024 30728
rect 7852 30688 8024 30716
rect 5074 30608 5080 30660
rect 5132 30608 5138 30660
rect 5813 30651 5871 30657
rect 5813 30617 5825 30651
rect 5859 30648 5871 30651
rect 6914 30648 6920 30660
rect 5859 30620 6920 30648
rect 5859 30617 5871 30620
rect 5813 30611 5871 30617
rect 6914 30608 6920 30620
rect 6972 30608 6978 30660
rect 7009 30651 7067 30657
rect 7009 30617 7021 30651
rect 7055 30648 7067 30651
rect 7098 30648 7104 30660
rect 7055 30620 7104 30648
rect 7055 30617 7067 30620
rect 7009 30611 7067 30617
rect 7098 30608 7104 30620
rect 7156 30608 7162 30660
rect 7282 30648 7288 30660
rect 7243 30620 7288 30648
rect 7282 30608 7288 30620
rect 7340 30648 7346 30660
rect 7852 30648 7880 30688
rect 8018 30676 8024 30688
rect 8076 30716 8082 30728
rect 8076 30688 8432 30716
rect 8076 30676 8082 30688
rect 7340 30620 7880 30648
rect 7340 30608 7346 30620
rect 7926 30608 7932 30660
rect 7984 30648 7990 30660
rect 8404 30657 8432 30688
rect 9766 30676 9772 30728
rect 9824 30716 9830 30728
rect 10873 30719 10931 30725
rect 10873 30716 10885 30719
rect 9824 30688 10885 30716
rect 9824 30676 9830 30688
rect 10873 30685 10885 30688
rect 10919 30685 10931 30719
rect 10873 30679 10931 30685
rect 11606 30676 11612 30728
rect 11664 30716 11670 30728
rect 11701 30719 11759 30725
rect 11701 30716 11713 30719
rect 11664 30688 11713 30716
rect 11664 30676 11670 30688
rect 11701 30685 11713 30688
rect 11747 30716 11759 30719
rect 11974 30716 11980 30728
rect 11747 30688 11980 30716
rect 11747 30685 11759 30688
rect 11701 30679 11759 30685
rect 11974 30676 11980 30688
rect 12032 30676 12038 30728
rect 8173 30651 8231 30657
rect 8173 30648 8185 30651
rect 7984 30620 8185 30648
rect 7984 30608 7990 30620
rect 8173 30617 8185 30620
rect 8219 30617 8231 30651
rect 8173 30611 8231 30617
rect 8389 30651 8447 30657
rect 8389 30617 8401 30651
rect 8435 30617 8447 30651
rect 9858 30648 9864 30660
rect 9819 30620 9864 30648
rect 8389 30611 8447 30617
rect 9858 30608 9864 30620
rect 9916 30608 9922 30660
rect 10597 30651 10655 30657
rect 10597 30617 10609 30651
rect 10643 30648 10655 30651
rect 12544 30648 12572 30824
rect 14090 30812 14096 30824
rect 14148 30812 14154 30864
rect 15746 30812 15752 30864
rect 15804 30852 15810 30864
rect 16209 30855 16267 30861
rect 16209 30852 16221 30855
rect 15804 30824 16221 30852
rect 15804 30812 15810 30824
rect 16209 30821 16221 30824
rect 16255 30852 16267 30855
rect 16255 30824 16344 30852
rect 16255 30821 16267 30824
rect 16209 30815 16267 30821
rect 12621 30787 12679 30793
rect 12621 30753 12633 30787
rect 12667 30784 12679 30787
rect 12710 30784 12716 30796
rect 12667 30756 12716 30784
rect 12667 30753 12679 30756
rect 12621 30747 12679 30753
rect 12710 30744 12716 30756
rect 12768 30744 12774 30796
rect 14182 30784 14188 30796
rect 12912 30756 14188 30784
rect 12802 30716 12808 30728
rect 12763 30688 12808 30716
rect 12802 30676 12808 30688
rect 12860 30676 12866 30728
rect 12912 30725 12940 30756
rect 14182 30744 14188 30756
rect 14240 30744 14246 30796
rect 16316 30784 16344 30824
rect 16666 30812 16672 30864
rect 16724 30852 16730 30864
rect 17589 30855 17647 30861
rect 17589 30852 17601 30855
rect 16724 30824 17601 30852
rect 16724 30812 16730 30824
rect 17589 30821 17601 30824
rect 17635 30852 17647 30855
rect 17862 30852 17868 30864
rect 17635 30824 17868 30852
rect 17635 30821 17647 30824
rect 17589 30815 17647 30821
rect 17862 30812 17868 30824
rect 17920 30812 17926 30864
rect 27080 30852 27108 30892
rect 29549 30889 29561 30923
rect 29595 30920 29607 30923
rect 30650 30920 30656 30932
rect 29595 30892 30656 30920
rect 29595 30889 29607 30892
rect 29549 30883 29607 30889
rect 30650 30880 30656 30892
rect 30708 30880 30714 30932
rect 36906 30920 36912 30932
rect 31726 30892 36912 30920
rect 31726 30852 31754 30892
rect 36906 30880 36912 30892
rect 36964 30880 36970 30932
rect 27080 30824 31754 30852
rect 18138 30784 18144 30796
rect 16316 30756 16896 30784
rect 18099 30756 18144 30784
rect 12897 30719 12955 30725
rect 12897 30685 12909 30719
rect 12943 30685 12955 30719
rect 12897 30679 12955 30685
rect 12986 30676 12992 30728
rect 13044 30716 13050 30728
rect 13265 30719 13323 30725
rect 13044 30688 13089 30716
rect 13044 30676 13050 30688
rect 13265 30685 13277 30719
rect 13311 30716 13323 30719
rect 13354 30716 13360 30728
rect 13311 30688 13360 30716
rect 13311 30685 13323 30688
rect 13265 30679 13323 30685
rect 13354 30676 13360 30688
rect 13412 30676 13418 30728
rect 14458 30716 14464 30728
rect 14419 30688 14464 30716
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 16868 30725 16896 30756
rect 18138 30744 18144 30756
rect 18196 30744 18202 30796
rect 18601 30787 18659 30793
rect 18601 30753 18613 30787
rect 18647 30784 18659 30787
rect 19150 30784 19156 30796
rect 18647 30756 19156 30784
rect 18647 30753 18659 30756
rect 18601 30747 18659 30753
rect 19150 30744 19156 30756
rect 19208 30744 19214 30796
rect 19242 30744 19248 30796
rect 19300 30784 19306 30796
rect 21453 30787 21511 30793
rect 21453 30784 21465 30787
rect 19300 30756 21465 30784
rect 19300 30744 19306 30756
rect 21453 30753 21465 30756
rect 21499 30753 21511 30787
rect 21453 30747 21511 30753
rect 26142 30744 26148 30796
rect 26200 30784 26206 30796
rect 27157 30787 27215 30793
rect 27157 30784 27169 30787
rect 26200 30756 27169 30784
rect 26200 30744 26206 30756
rect 27157 30753 27169 30756
rect 27203 30753 27215 30787
rect 27157 30747 27215 30753
rect 28350 30744 28356 30796
rect 28408 30784 28414 30796
rect 28629 30787 28687 30793
rect 28629 30784 28641 30787
rect 28408 30756 28641 30784
rect 28408 30744 28414 30756
rect 28629 30753 28641 30756
rect 28675 30753 28687 30787
rect 33410 30784 33416 30796
rect 28629 30747 28687 30753
rect 29656 30756 30144 30784
rect 16853 30719 16911 30725
rect 16853 30685 16865 30719
rect 16899 30685 16911 30719
rect 16853 30679 16911 30685
rect 17034 30676 17040 30728
rect 17092 30716 17098 30728
rect 17405 30719 17463 30725
rect 17405 30716 17417 30719
rect 17092 30688 17417 30716
rect 17092 30676 17098 30688
rect 17405 30685 17417 30688
rect 17451 30716 17463 30719
rect 17586 30716 17592 30728
rect 17451 30688 17592 30716
rect 17451 30685 17463 30688
rect 17405 30679 17463 30685
rect 17586 30676 17592 30688
rect 17644 30676 17650 30728
rect 18046 30676 18052 30728
rect 18104 30716 18110 30728
rect 18233 30719 18291 30725
rect 18233 30716 18245 30719
rect 18104 30688 18245 30716
rect 18104 30676 18110 30688
rect 18233 30685 18245 30688
rect 18279 30716 18291 30719
rect 19260 30716 19288 30744
rect 18279 30688 19288 30716
rect 18279 30685 18291 30688
rect 18233 30679 18291 30685
rect 19426 30676 19432 30728
rect 19484 30716 19490 30728
rect 19705 30719 19763 30725
rect 19705 30716 19717 30719
rect 19484 30688 19717 30716
rect 19484 30676 19490 30688
rect 19705 30685 19717 30688
rect 19751 30685 19763 30719
rect 21913 30719 21971 30725
rect 21913 30716 21925 30719
rect 19705 30679 19763 30685
rect 21284 30688 21925 30716
rect 13107 30651 13165 30657
rect 13107 30648 13119 30651
rect 10643 30620 12572 30648
rect 12728 30620 13119 30648
rect 10643 30617 10655 30620
rect 10597 30611 10655 30617
rect 4341 30583 4399 30589
rect 4341 30549 4353 30583
rect 4387 30580 4399 30583
rect 5902 30580 5908 30592
rect 4387 30552 5908 30580
rect 4387 30549 4399 30552
rect 4341 30543 4399 30549
rect 5902 30540 5908 30552
rect 5960 30540 5966 30592
rect 7374 30580 7380 30592
rect 7335 30552 7380 30580
rect 7374 30540 7380 30552
rect 7432 30540 7438 30592
rect 7834 30540 7840 30592
rect 7892 30580 7898 30592
rect 8021 30583 8079 30589
rect 8021 30580 8033 30583
rect 7892 30552 8033 30580
rect 7892 30540 7898 30552
rect 8021 30549 8033 30552
rect 8067 30549 8079 30583
rect 8021 30543 8079 30549
rect 9661 30583 9719 30589
rect 9661 30549 9673 30583
rect 9707 30580 9719 30583
rect 10410 30580 10416 30592
rect 9707 30552 10416 30580
rect 9707 30549 9719 30552
rect 9661 30543 9719 30549
rect 10410 30540 10416 30552
rect 10468 30540 10474 30592
rect 11882 30580 11888 30592
rect 11843 30552 11888 30580
rect 11882 30540 11888 30552
rect 11940 30540 11946 30592
rect 12066 30540 12072 30592
rect 12124 30580 12130 30592
rect 12250 30580 12256 30592
rect 12124 30552 12256 30580
rect 12124 30540 12130 30552
rect 12250 30540 12256 30552
rect 12308 30580 12314 30592
rect 12728 30580 12756 30620
rect 13107 30617 13119 30620
rect 13153 30617 13165 30651
rect 14734 30648 14740 30660
rect 14695 30620 14740 30648
rect 13107 30611 13165 30617
rect 14734 30608 14740 30620
rect 14792 30608 14798 30660
rect 17126 30648 17132 30660
rect 15962 30620 17132 30648
rect 17126 30608 17132 30620
rect 17184 30608 17190 30660
rect 19978 30648 19984 30660
rect 19939 30620 19984 30648
rect 19978 30608 19984 30620
rect 20036 30608 20042 30660
rect 20990 30608 20996 30660
rect 21048 30608 21054 30660
rect 12308 30552 12756 30580
rect 12308 30540 12314 30552
rect 15010 30540 15016 30592
rect 15068 30580 15074 30592
rect 16669 30583 16727 30589
rect 16669 30580 16681 30583
rect 15068 30552 16681 30580
rect 15068 30540 15074 30552
rect 16669 30549 16681 30552
rect 16715 30549 16727 30583
rect 16669 30543 16727 30549
rect 20806 30540 20812 30592
rect 20864 30580 20870 30592
rect 21284 30580 21312 30688
rect 21913 30685 21925 30688
rect 21959 30685 21971 30719
rect 21913 30679 21971 30685
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30716 24823 30719
rect 25130 30716 25136 30728
rect 24811 30688 25136 30716
rect 24811 30685 24823 30688
rect 24765 30679 24823 30685
rect 25130 30676 25136 30688
rect 25188 30676 25194 30728
rect 28445 30719 28503 30725
rect 28445 30685 28457 30719
rect 28491 30716 28503 30719
rect 29178 30716 29184 30728
rect 28491 30688 29184 30716
rect 28491 30685 28503 30688
rect 28445 30679 28503 30685
rect 29178 30676 29184 30688
rect 29236 30676 29242 30728
rect 22186 30648 22192 30660
rect 22147 30620 22192 30648
rect 22186 30608 22192 30620
rect 22244 30608 22250 30660
rect 22922 30608 22928 30660
rect 22980 30608 22986 30660
rect 24946 30608 24952 30660
rect 25004 30648 25010 30660
rect 26881 30651 26939 30657
rect 25004 30620 25714 30648
rect 25004 30608 25010 30620
rect 26881 30617 26893 30651
rect 26927 30648 26939 30651
rect 27982 30648 27988 30660
rect 26927 30620 27988 30648
rect 26927 30617 26939 30620
rect 26881 30611 26939 30617
rect 27982 30608 27988 30620
rect 28040 30608 28046 30660
rect 28353 30651 28411 30657
rect 28353 30617 28365 30651
rect 28399 30648 28411 30651
rect 28902 30648 28908 30660
rect 28399 30620 28908 30648
rect 28399 30617 28411 30620
rect 28353 30611 28411 30617
rect 28902 30608 28908 30620
rect 28960 30648 28966 30660
rect 29656 30648 29684 30756
rect 29733 30719 29791 30725
rect 29733 30685 29745 30719
rect 29779 30685 29791 30719
rect 29914 30716 29920 30728
rect 29875 30688 29920 30716
rect 29733 30679 29791 30685
rect 28960 30620 29684 30648
rect 28960 30608 28966 30620
rect 20864 30552 21312 30580
rect 24857 30583 24915 30589
rect 20864 30540 20870 30552
rect 24857 30549 24869 30583
rect 24903 30580 24915 30583
rect 25314 30580 25320 30592
rect 24903 30552 25320 30580
rect 24903 30549 24915 30552
rect 24857 30543 24915 30549
rect 25314 30540 25320 30552
rect 25372 30540 25378 30592
rect 25409 30583 25467 30589
rect 25409 30549 25421 30583
rect 25455 30580 25467 30583
rect 26786 30580 26792 30592
rect 25455 30552 26792 30580
rect 25455 30549 25467 30552
rect 25409 30543 25467 30549
rect 26786 30540 26792 30552
rect 26844 30540 26850 30592
rect 27062 30540 27068 30592
rect 27120 30580 27126 30592
rect 28077 30583 28135 30589
rect 28077 30580 28089 30583
rect 27120 30552 28089 30580
rect 27120 30540 27126 30552
rect 28077 30549 28089 30552
rect 28123 30549 28135 30583
rect 28258 30580 28264 30592
rect 28219 30552 28264 30580
rect 28077 30543 28135 30549
rect 28258 30540 28264 30552
rect 28316 30540 28322 30592
rect 29748 30580 29776 30679
rect 29914 30676 29920 30688
rect 29972 30676 29978 30728
rect 30116 30725 30144 30756
rect 31726 30756 33416 30784
rect 30101 30719 30159 30725
rect 30101 30685 30113 30719
rect 30147 30716 30159 30719
rect 30190 30716 30196 30728
rect 30147 30688 30196 30716
rect 30147 30685 30159 30688
rect 30101 30679 30159 30685
rect 30190 30676 30196 30688
rect 30248 30676 30254 30728
rect 30374 30676 30380 30728
rect 30432 30716 30438 30728
rect 30926 30716 30932 30728
rect 30432 30688 30932 30716
rect 30432 30676 30438 30688
rect 30926 30676 30932 30688
rect 30984 30716 30990 30728
rect 31297 30719 31355 30725
rect 31297 30716 31309 30719
rect 30984 30688 31309 30716
rect 30984 30676 30990 30688
rect 31297 30685 31309 30688
rect 31343 30716 31355 30719
rect 31726 30716 31754 30756
rect 33410 30744 33416 30756
rect 33468 30784 33474 30796
rect 33468 30756 33824 30784
rect 33468 30744 33474 30756
rect 33796 30725 33824 30756
rect 35434 30744 35440 30796
rect 35492 30784 35498 30796
rect 36265 30787 36323 30793
rect 36265 30784 36277 30787
rect 35492 30756 36277 30784
rect 35492 30744 35498 30756
rect 36265 30753 36277 30756
rect 36311 30753 36323 30787
rect 36446 30784 36452 30796
rect 36407 30756 36452 30784
rect 36265 30747 36323 30753
rect 36446 30744 36452 30756
rect 36504 30744 36510 30796
rect 31343 30688 31754 30716
rect 33781 30719 33839 30725
rect 31343 30685 31355 30688
rect 31297 30679 31355 30685
rect 33781 30685 33793 30719
rect 33827 30716 33839 30719
rect 34238 30716 34244 30728
rect 33827 30688 34244 30716
rect 33827 30685 33839 30688
rect 33781 30679 33839 30685
rect 34238 30676 34244 30688
rect 34296 30676 34302 30728
rect 34606 30676 34612 30728
rect 34664 30716 34670 30728
rect 35253 30719 35311 30725
rect 35253 30716 35265 30719
rect 34664 30688 35265 30716
rect 34664 30676 34670 30688
rect 35253 30685 35265 30688
rect 35299 30716 35311 30719
rect 35526 30716 35532 30728
rect 35299 30688 35532 30716
rect 35299 30685 35311 30688
rect 35253 30679 35311 30685
rect 35526 30676 35532 30688
rect 35584 30676 35590 30728
rect 29822 30608 29828 30660
rect 29880 30648 29886 30660
rect 29880 30620 29925 30648
rect 29880 30608 29886 30620
rect 30282 30608 30288 30660
rect 30340 30648 30346 30660
rect 30561 30651 30619 30657
rect 30561 30648 30573 30651
rect 30340 30620 30573 30648
rect 30340 30608 30346 30620
rect 30561 30617 30573 30620
rect 30607 30617 30619 30651
rect 30742 30648 30748 30660
rect 30703 30620 30748 30648
rect 30561 30611 30619 30617
rect 30742 30608 30748 30620
rect 30800 30608 30806 30660
rect 31481 30651 31539 30657
rect 31481 30617 31493 30651
rect 31527 30648 31539 30651
rect 32214 30648 32220 30660
rect 31527 30620 32220 30648
rect 31527 30617 31539 30620
rect 31481 30611 31539 30617
rect 32214 30608 32220 30620
rect 32272 30608 32278 30660
rect 33042 30608 33048 30660
rect 33100 30608 33106 30660
rect 33502 30648 33508 30660
rect 33463 30620 33508 30648
rect 33502 30608 33508 30620
rect 33560 30608 33566 30660
rect 38102 30648 38108 30660
rect 38063 30620 38108 30648
rect 38102 30608 38108 30620
rect 38160 30608 38166 30660
rect 30466 30580 30472 30592
rect 29748 30552 30472 30580
rect 30466 30540 30472 30552
rect 30524 30540 30530 30592
rect 32030 30580 32036 30592
rect 31991 30552 32036 30580
rect 32030 30540 32036 30552
rect 32088 30540 32094 30592
rect 35250 30540 35256 30592
rect 35308 30580 35314 30592
rect 35345 30583 35403 30589
rect 35345 30580 35357 30583
rect 35308 30552 35357 30580
rect 35308 30540 35314 30552
rect 35345 30549 35357 30552
rect 35391 30549 35403 30583
rect 35345 30543 35403 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 6914 30336 6920 30388
rect 6972 30376 6978 30388
rect 7837 30379 7895 30385
rect 7837 30376 7849 30379
rect 6972 30348 7849 30376
rect 6972 30336 6978 30348
rect 7837 30345 7849 30348
rect 7883 30345 7895 30379
rect 7837 30339 7895 30345
rect 8018 30336 8024 30388
rect 8076 30336 8082 30388
rect 10413 30379 10471 30385
rect 10413 30345 10425 30379
rect 10459 30376 10471 30379
rect 10594 30376 10600 30388
rect 10459 30348 10600 30376
rect 10459 30345 10471 30348
rect 10413 30339 10471 30345
rect 10594 30336 10600 30348
rect 10652 30336 10658 30388
rect 12802 30376 12808 30388
rect 12763 30348 12808 30376
rect 12802 30336 12808 30348
rect 12860 30336 12866 30388
rect 14182 30336 14188 30388
rect 14240 30376 14246 30388
rect 14277 30379 14335 30385
rect 14277 30376 14289 30379
rect 14240 30348 14289 30376
rect 14240 30336 14246 30348
rect 14277 30345 14289 30348
rect 14323 30345 14335 30379
rect 14277 30339 14335 30345
rect 14734 30336 14740 30388
rect 14792 30376 14798 30388
rect 14921 30379 14979 30385
rect 14921 30376 14933 30379
rect 14792 30348 14933 30376
rect 14792 30336 14798 30348
rect 14921 30345 14933 30348
rect 14967 30345 14979 30379
rect 14921 30339 14979 30345
rect 15028 30348 15608 30376
rect 5353 30311 5411 30317
rect 5353 30277 5365 30311
rect 5399 30308 5411 30311
rect 7374 30308 7380 30320
rect 5399 30280 7380 30308
rect 5399 30277 5411 30280
rect 5353 30271 5411 30277
rect 7374 30268 7380 30280
rect 7432 30268 7438 30320
rect 8036 30308 8064 30336
rect 8113 30311 8171 30317
rect 8113 30308 8125 30311
rect 8036 30280 8125 30308
rect 8113 30277 8125 30280
rect 8159 30277 8171 30311
rect 8113 30271 8171 30277
rect 12158 30268 12164 30320
rect 12216 30308 12222 30320
rect 13262 30308 13268 30320
rect 12216 30280 12664 30308
rect 13223 30280 13268 30308
rect 12216 30268 12222 30280
rect 4893 30243 4951 30249
rect 4893 30209 4905 30243
rect 4939 30240 4951 30243
rect 5166 30240 5172 30252
rect 4939 30212 5172 30240
rect 4939 30209 4951 30212
rect 4893 30203 4951 30209
rect 5166 30200 5172 30212
rect 5224 30200 5230 30252
rect 5629 30243 5687 30249
rect 5629 30209 5641 30243
rect 5675 30240 5687 30243
rect 6825 30243 6883 30249
rect 5675 30212 6684 30240
rect 5675 30209 5687 30212
rect 5629 30203 5687 30209
rect 5537 30175 5595 30181
rect 5537 30141 5549 30175
rect 5583 30172 5595 30175
rect 5902 30172 5908 30184
rect 5583 30144 5908 30172
rect 5583 30141 5595 30144
rect 5537 30135 5595 30141
rect 5902 30132 5908 30144
rect 5960 30132 5966 30184
rect 6549 30175 6607 30181
rect 6549 30141 6561 30175
rect 6595 30141 6607 30175
rect 6656 30172 6684 30212
rect 6825 30209 6837 30243
rect 6871 30240 6883 30243
rect 7466 30240 7472 30252
rect 6871 30212 7472 30240
rect 6871 30209 6883 30212
rect 6825 30203 6883 30209
rect 7466 30200 7472 30212
rect 7524 30200 7530 30252
rect 8021 30243 8079 30249
rect 8021 30240 8033 30243
rect 7944 30212 8033 30240
rect 7098 30172 7104 30184
rect 6656 30144 7104 30172
rect 6549 30135 6607 30141
rect 6564 30104 6592 30135
rect 7098 30132 7104 30144
rect 7156 30132 7162 30184
rect 5644 30076 6592 30104
rect 4798 30036 4804 30048
rect 4759 30008 4804 30036
rect 4798 29996 4804 30008
rect 4856 29996 4862 30048
rect 4890 29996 4896 30048
rect 4948 30036 4954 30048
rect 5644 30045 5672 30076
rect 7006 30064 7012 30116
rect 7064 30104 7070 30116
rect 7944 30104 7972 30212
rect 8021 30209 8033 30212
rect 8067 30209 8079 30243
rect 8021 30203 8079 30209
rect 8205 30243 8263 30249
rect 8205 30209 8217 30243
rect 8251 30209 8263 30243
rect 8386 30240 8392 30252
rect 8347 30212 8392 30240
rect 8205 30203 8263 30209
rect 8220 30172 8248 30203
rect 8386 30200 8392 30212
rect 8444 30200 8450 30252
rect 9674 30200 9680 30252
rect 9732 30240 9738 30252
rect 9858 30240 9864 30252
rect 9732 30212 9864 30240
rect 9732 30200 9738 30212
rect 9858 30200 9864 30212
rect 9916 30240 9922 30252
rect 9953 30243 10011 30249
rect 9953 30240 9965 30243
rect 9916 30212 9965 30240
rect 9916 30200 9922 30212
rect 9953 30209 9965 30212
rect 9999 30209 10011 30243
rect 10226 30240 10232 30252
rect 10187 30212 10232 30240
rect 9953 30203 10011 30209
rect 10226 30200 10232 30212
rect 10284 30200 10290 30252
rect 11514 30240 11520 30252
rect 11475 30212 11520 30240
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 11609 30243 11667 30249
rect 11609 30209 11621 30243
rect 11655 30240 11667 30243
rect 11882 30240 11888 30252
rect 11655 30212 11888 30240
rect 11655 30209 11667 30212
rect 11609 30203 11667 30209
rect 11882 30200 11888 30212
rect 11940 30200 11946 30252
rect 12342 30240 12348 30252
rect 12303 30212 12348 30240
rect 12342 30200 12348 30212
rect 12400 30200 12406 30252
rect 12636 30249 12664 30280
rect 13262 30268 13268 30280
rect 13320 30268 13326 30320
rect 13446 30308 13452 30320
rect 13504 30317 13510 30320
rect 13504 30311 13539 30317
rect 13391 30280 13452 30308
rect 13446 30268 13452 30280
rect 13527 30308 13539 30311
rect 15028 30308 15056 30348
rect 15194 30308 15200 30320
rect 13527 30280 15056 30308
rect 15155 30280 15200 30308
rect 13527 30277 13539 30280
rect 13504 30271 13539 30277
rect 13504 30268 13510 30271
rect 15194 30268 15200 30280
rect 15252 30268 15258 30320
rect 15378 30268 15384 30320
rect 15436 30317 15442 30320
rect 15436 30311 15465 30317
rect 15453 30277 15465 30311
rect 15436 30271 15465 30277
rect 15436 30268 15442 30271
rect 12620 30243 12678 30249
rect 12620 30209 12632 30243
rect 12666 30209 12678 30243
rect 12620 30203 12678 30209
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 14185 30243 14243 30249
rect 14185 30240 14197 30243
rect 14056 30212 14197 30240
rect 14056 30200 14062 30212
rect 14185 30209 14197 30212
rect 14231 30209 14243 30243
rect 14185 30203 14243 30209
rect 14461 30243 14519 30249
rect 14461 30209 14473 30243
rect 14507 30240 14519 30243
rect 14734 30240 14740 30252
rect 14507 30212 14740 30240
rect 14507 30209 14519 30212
rect 14461 30203 14519 30209
rect 14734 30200 14740 30212
rect 14792 30200 14798 30252
rect 15105 30243 15163 30249
rect 15105 30209 15117 30243
rect 15151 30209 15163 30243
rect 15286 30240 15292 30252
rect 15247 30212 15292 30240
rect 15105 30203 15163 30209
rect 10042 30172 10048 30184
rect 8036 30144 8248 30172
rect 10003 30144 10048 30172
rect 8036 30116 8064 30144
rect 10042 30132 10048 30144
rect 10100 30132 10106 30184
rect 11146 30132 11152 30184
rect 11204 30172 11210 30184
rect 11793 30175 11851 30181
rect 11793 30172 11805 30175
rect 11204 30144 11805 30172
rect 11204 30132 11210 30144
rect 11793 30141 11805 30144
rect 11839 30141 11851 30175
rect 11793 30135 11851 30141
rect 7064 30076 7972 30104
rect 7064 30064 7070 30076
rect 8018 30064 8024 30116
rect 8076 30064 8082 30116
rect 11422 30064 11428 30116
rect 11480 30104 11486 30116
rect 11606 30104 11612 30116
rect 11480 30076 11612 30104
rect 11480 30064 11486 30076
rect 11606 30064 11612 30076
rect 11664 30064 11670 30116
rect 11808 30104 11836 30135
rect 12250 30132 12256 30184
rect 12308 30172 12314 30184
rect 12436 30175 12494 30181
rect 12308 30164 12388 30172
rect 12436 30164 12448 30175
rect 12308 30144 12448 30164
rect 12308 30132 12314 30144
rect 12360 30141 12448 30144
rect 12482 30141 12494 30175
rect 12360 30136 12494 30141
rect 12436 30135 12494 30136
rect 12526 30132 12532 30184
rect 12584 30172 12590 30184
rect 15120 30172 15148 30203
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 15580 30240 15608 30348
rect 19426 30336 19432 30388
rect 19484 30336 19490 30388
rect 19705 30379 19763 30385
rect 19705 30345 19717 30379
rect 19751 30376 19763 30379
rect 19978 30376 19984 30388
rect 19751 30348 19984 30376
rect 19751 30345 19763 30348
rect 19705 30339 19763 30345
rect 19978 30336 19984 30348
rect 20036 30336 20042 30388
rect 20990 30376 20996 30388
rect 20916 30348 20996 30376
rect 16482 30268 16488 30320
rect 16540 30308 16546 30320
rect 17037 30311 17095 30317
rect 17037 30308 17049 30311
rect 16540 30280 17049 30308
rect 16540 30268 16546 30280
rect 17037 30277 17049 30280
rect 17083 30277 17095 30311
rect 17037 30271 17095 30277
rect 17310 30268 17316 30320
rect 17368 30308 17374 30320
rect 19444 30308 19472 30336
rect 20806 30308 20812 30320
rect 17368 30280 20812 30308
rect 17368 30268 17374 30280
rect 20806 30268 20812 30280
rect 20864 30268 20870 30320
rect 20916 30317 20944 30348
rect 20990 30336 20996 30348
rect 21048 30336 21054 30388
rect 22186 30336 22192 30388
rect 22244 30376 22250 30388
rect 22373 30379 22431 30385
rect 22373 30376 22385 30379
rect 22244 30348 22385 30376
rect 22244 30336 22250 30348
rect 22373 30345 22385 30348
rect 22419 30345 22431 30379
rect 27154 30376 27160 30388
rect 22373 30339 22431 30345
rect 27080 30348 27160 30376
rect 20901 30311 20959 30317
rect 20901 30277 20913 30311
rect 20947 30277 20959 30311
rect 20901 30271 20959 30277
rect 22922 30268 22928 30320
rect 22980 30308 22986 30320
rect 23109 30311 23167 30317
rect 23109 30308 23121 30311
rect 22980 30280 23121 30308
rect 22980 30268 22986 30280
rect 23109 30277 23121 30280
rect 23155 30277 23167 30311
rect 23109 30271 23167 30277
rect 25961 30311 26019 30317
rect 25961 30277 25973 30311
rect 26007 30308 26019 30311
rect 26973 30311 27031 30317
rect 26973 30308 26985 30311
rect 26007 30280 26985 30308
rect 26007 30277 26019 30280
rect 25961 30271 26019 30277
rect 26973 30277 26985 30280
rect 27019 30277 27031 30311
rect 26973 30271 27031 30277
rect 27080 30262 27108 30348
rect 27154 30336 27160 30348
rect 27212 30336 27218 30388
rect 29178 30336 29184 30388
rect 29236 30376 29242 30388
rect 30006 30376 30012 30388
rect 29236 30348 30012 30376
rect 29236 30336 29242 30348
rect 30006 30336 30012 30348
rect 30064 30336 30070 30388
rect 30282 30336 30288 30388
rect 30340 30376 30346 30388
rect 30340 30348 31432 30376
rect 30340 30336 30346 30348
rect 27158 30265 27216 30271
rect 27246 30268 27252 30320
rect 27304 30308 27310 30320
rect 27304 30280 27349 30308
rect 27304 30268 27310 30280
rect 27430 30268 27436 30320
rect 27488 30317 27494 30320
rect 27488 30311 27517 30317
rect 27505 30277 27517 30311
rect 27488 30271 27517 30277
rect 27488 30268 27494 30271
rect 27706 30268 27712 30320
rect 27764 30308 27770 30320
rect 28169 30311 28227 30317
rect 28169 30308 28181 30311
rect 27764 30280 28181 30308
rect 27764 30268 27770 30280
rect 28169 30277 28181 30280
rect 28215 30277 28227 30311
rect 28994 30308 29000 30320
rect 28955 30280 29000 30308
rect 28169 30271 28227 30277
rect 28994 30268 29000 30280
rect 29052 30268 29058 30320
rect 30374 30308 30380 30320
rect 29840 30280 30380 30308
rect 27158 30262 27170 30265
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 15580 30212 16957 30240
rect 16945 30209 16957 30212
rect 16991 30209 17003 30243
rect 16945 30203 17003 30209
rect 17129 30243 17187 30249
rect 17129 30209 17141 30243
rect 17175 30240 17187 30243
rect 18046 30240 18052 30252
rect 17175 30212 18052 30240
rect 17175 30209 17187 30212
rect 17129 30203 17187 30209
rect 18046 30200 18052 30212
rect 18104 30200 18110 30252
rect 18414 30240 18420 30252
rect 18375 30212 18420 30240
rect 18414 30200 18420 30212
rect 18472 30200 18478 30252
rect 18598 30200 18604 30252
rect 18656 30240 18662 30252
rect 18693 30243 18751 30249
rect 18693 30240 18705 30243
rect 18656 30212 18705 30240
rect 18656 30200 18662 30212
rect 18693 30209 18705 30212
rect 18739 30209 18751 30243
rect 19150 30240 19156 30252
rect 19111 30212 19156 30240
rect 18693 30203 18751 30209
rect 19150 30200 19156 30212
rect 19208 30200 19214 30252
rect 19334 30240 19340 30252
rect 19295 30212 19340 30240
rect 19334 30200 19340 30212
rect 19392 30200 19398 30252
rect 19429 30243 19487 30249
rect 19429 30209 19441 30243
rect 19475 30209 19487 30243
rect 19429 30203 19487 30209
rect 19521 30243 19579 30249
rect 19521 30209 19533 30243
rect 19567 30240 19579 30243
rect 19610 30240 19616 30252
rect 19567 30212 19616 30240
rect 19567 30209 19579 30212
rect 19521 30203 19579 30209
rect 15470 30172 15476 30184
rect 12584 30144 12628 30172
rect 15120 30144 15476 30172
rect 12584 30132 12590 30144
rect 15470 30132 15476 30144
rect 15528 30132 15534 30184
rect 15565 30175 15623 30181
rect 15565 30141 15577 30175
rect 15611 30172 15623 30175
rect 15654 30172 15660 30184
rect 15611 30144 15660 30172
rect 15611 30141 15623 30144
rect 15565 30135 15623 30141
rect 15654 30132 15660 30144
rect 15712 30132 15718 30184
rect 16758 30172 16764 30184
rect 16719 30144 16764 30172
rect 16758 30132 16764 30144
rect 16816 30132 16822 30184
rect 17313 30175 17371 30181
rect 17313 30141 17325 30175
rect 17359 30172 17371 30175
rect 18138 30172 18144 30184
rect 17359 30144 18144 30172
rect 17359 30141 17371 30144
rect 17313 30135 17371 30141
rect 18138 30132 18144 30144
rect 18196 30132 18202 30184
rect 18506 30172 18512 30184
rect 18467 30144 18512 30172
rect 18506 30132 18512 30144
rect 18564 30132 18570 30184
rect 19242 30132 19248 30184
rect 19300 30172 19306 30184
rect 19444 30172 19472 30203
rect 19610 30200 19616 30212
rect 19668 30240 19674 30252
rect 20070 30240 20076 30252
rect 19668 30212 20076 30240
rect 19668 30200 19674 30212
rect 20070 30200 20076 30212
rect 20128 30200 20134 30252
rect 20162 30200 20168 30252
rect 20220 30240 20226 30252
rect 20220 30212 20265 30240
rect 20220 30200 20226 30212
rect 20714 30200 20720 30252
rect 20772 30240 20778 30252
rect 20993 30243 21051 30249
rect 20993 30240 21005 30243
rect 20772 30212 21005 30240
rect 20772 30200 20778 30212
rect 20993 30209 21005 30212
rect 21039 30240 21051 30243
rect 22554 30240 22560 30252
rect 21039 30212 22094 30240
rect 22515 30212 22560 30240
rect 21039 30209 21051 30212
rect 20993 30203 21051 30209
rect 19300 30144 19472 30172
rect 22066 30172 22094 30212
rect 22554 30200 22560 30212
rect 22612 30200 22618 30252
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30240 23259 30243
rect 23382 30240 23388 30252
rect 23247 30212 23388 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 23382 30200 23388 30212
rect 23440 30240 23446 30252
rect 23845 30243 23903 30249
rect 23845 30240 23857 30243
rect 23440 30212 23857 30240
rect 23440 30200 23446 30212
rect 23845 30209 23857 30212
rect 23891 30209 23903 30243
rect 23845 30203 23903 30209
rect 24854 30200 24860 30252
rect 24912 30200 24918 30252
rect 27080 30234 27170 30262
rect 27158 30231 27170 30234
rect 27204 30231 27216 30265
rect 27158 30225 27216 30231
rect 27341 30243 27399 30249
rect 27341 30209 27353 30243
rect 27387 30230 27399 30243
rect 28074 30240 28080 30252
rect 27387 30209 27416 30230
rect 28035 30212 28080 30240
rect 27341 30203 27416 30209
rect 27356 30202 27416 30203
rect 22830 30172 22836 30184
rect 22066 30144 22836 30172
rect 19300 30132 19306 30144
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 23937 30175 23995 30181
rect 23937 30141 23949 30175
rect 23983 30172 23995 30175
rect 24946 30172 24952 30184
rect 23983 30144 24952 30172
rect 23983 30141 23995 30144
rect 23937 30135 23995 30141
rect 24946 30132 24952 30144
rect 25004 30132 25010 30184
rect 26234 30172 26240 30184
rect 26195 30144 26240 30172
rect 26234 30132 26240 30144
rect 26292 30132 26298 30184
rect 18230 30104 18236 30116
rect 11808 30076 14964 30104
rect 18191 30076 18236 30104
rect 5629 30039 5687 30045
rect 5629 30036 5641 30039
rect 4948 30008 5641 30036
rect 4948 29996 4954 30008
rect 5629 30005 5641 30008
rect 5675 30005 5687 30039
rect 5629 29999 5687 30005
rect 5813 30039 5871 30045
rect 5813 30005 5825 30039
rect 5859 30036 5871 30039
rect 9766 30036 9772 30048
rect 5859 30008 9772 30036
rect 5859 30005 5871 30008
rect 5813 29999 5871 30005
rect 9766 29996 9772 30008
rect 9824 29996 9830 30048
rect 10229 30039 10287 30045
rect 10229 30005 10241 30039
rect 10275 30036 10287 30039
rect 11514 30036 11520 30048
rect 10275 30008 11520 30036
rect 10275 30005 10287 30008
rect 10229 29999 10287 30005
rect 11514 29996 11520 30008
rect 11572 29996 11578 30048
rect 11701 30039 11759 30045
rect 11701 30005 11713 30039
rect 11747 30036 11759 30039
rect 11790 30036 11796 30048
rect 11747 30008 11796 30036
rect 11747 30005 11759 30008
rect 11701 29999 11759 30005
rect 11790 29996 11796 30008
rect 11848 29996 11854 30048
rect 11974 29996 11980 30048
rect 12032 30036 12038 30048
rect 13449 30039 13507 30045
rect 13449 30036 13461 30039
rect 12032 30008 13461 30036
rect 12032 29996 12038 30008
rect 13449 30005 13461 30008
rect 13495 30005 13507 30039
rect 13630 30036 13636 30048
rect 13591 30008 13636 30036
rect 13449 29999 13507 30005
rect 13630 29996 13636 30008
rect 13688 29996 13694 30048
rect 13814 29996 13820 30048
rect 13872 30036 13878 30048
rect 14461 30039 14519 30045
rect 14461 30036 14473 30039
rect 13872 30008 14473 30036
rect 13872 29996 13878 30008
rect 14461 30005 14473 30008
rect 14507 30005 14519 30039
rect 14936 30036 14964 30076
rect 18230 30064 18236 30076
rect 18288 30064 18294 30116
rect 20257 30107 20315 30113
rect 20257 30104 20269 30107
rect 18340 30076 20269 30104
rect 17034 30036 17040 30048
rect 14936 30008 17040 30036
rect 14461 29999 14519 30005
rect 17034 29996 17040 30008
rect 17092 29996 17098 30048
rect 17126 29996 17132 30048
rect 17184 30036 17190 30048
rect 18340 30036 18368 30076
rect 20257 30073 20269 30076
rect 20303 30073 20315 30107
rect 20257 30067 20315 30073
rect 26418 30064 26424 30116
rect 26476 30104 26482 30116
rect 27388 30104 27416 30202
rect 28074 30200 28080 30212
rect 28132 30200 28138 30252
rect 29840 30249 29868 30280
rect 30374 30268 30380 30280
rect 30432 30268 30438 30320
rect 30834 30268 30840 30320
rect 30892 30268 30898 30320
rect 28905 30243 28963 30249
rect 28905 30209 28917 30243
rect 28951 30209 28963 30243
rect 28905 30203 28963 30209
rect 29089 30243 29147 30249
rect 29089 30209 29101 30243
rect 29135 30209 29147 30243
rect 29089 30203 29147 30209
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 31404 30240 31432 30348
rect 31846 30336 31852 30388
rect 31904 30376 31910 30388
rect 32582 30376 32588 30388
rect 31904 30348 32588 30376
rect 31904 30336 31910 30348
rect 32582 30336 32588 30348
rect 32640 30336 32646 30388
rect 35526 30336 35532 30388
rect 35584 30376 35590 30388
rect 35584 30348 35848 30376
rect 35584 30336 35590 30348
rect 31478 30268 31484 30320
rect 31536 30308 31542 30320
rect 33781 30311 33839 30317
rect 31536 30280 33640 30308
rect 31536 30268 31542 30280
rect 33612 30249 33640 30280
rect 33781 30277 33793 30311
rect 33827 30308 33839 30311
rect 34517 30311 34575 30317
rect 34517 30308 34529 30311
rect 33827 30280 34529 30308
rect 33827 30277 33839 30280
rect 33781 30271 33839 30277
rect 34517 30277 34529 30280
rect 34563 30277 34575 30311
rect 34517 30271 34575 30277
rect 35250 30268 35256 30320
rect 35308 30268 35314 30320
rect 32217 30243 32275 30249
rect 32217 30240 32229 30243
rect 31404 30212 32229 30240
rect 29825 30203 29883 30209
rect 32217 30209 32229 30212
rect 32263 30209 32275 30243
rect 32217 30203 32275 30209
rect 33597 30243 33655 30249
rect 33597 30209 33609 30243
rect 33643 30209 33655 30243
rect 35820 30240 35848 30348
rect 36449 30243 36507 30249
rect 36449 30240 36461 30243
rect 35820 30212 36461 30240
rect 33597 30203 33655 30209
rect 36449 30209 36461 30212
rect 36495 30209 36507 30243
rect 37550 30240 37556 30252
rect 37511 30212 37556 30240
rect 36449 30203 36507 30209
rect 27617 30175 27675 30181
rect 27617 30141 27629 30175
rect 27663 30141 27675 30175
rect 28920 30172 28948 30203
rect 28920 30144 29040 30172
rect 27617 30135 27675 30141
rect 26476 30076 27416 30104
rect 27632 30104 27660 30135
rect 29012 30116 29040 30144
rect 27890 30104 27896 30116
rect 27632 30076 27896 30104
rect 26476 30064 26482 30076
rect 27890 30064 27896 30076
rect 27948 30064 27954 30116
rect 28994 30064 29000 30116
rect 29052 30064 29058 30116
rect 17184 30008 18368 30036
rect 18693 30039 18751 30045
rect 17184 29996 17190 30008
rect 18693 30005 18705 30039
rect 18739 30036 18751 30039
rect 19242 30036 19248 30048
rect 18739 30008 19248 30036
rect 18739 30005 18751 30008
rect 18693 29999 18751 30005
rect 19242 29996 19248 30008
rect 19300 29996 19306 30048
rect 24489 30039 24547 30045
rect 24489 30005 24501 30039
rect 24535 30036 24547 30039
rect 26602 30036 26608 30048
rect 24535 30008 26608 30036
rect 24535 30005 24547 30008
rect 24489 29999 24547 30005
rect 26602 29996 26608 30008
rect 26660 30036 26666 30048
rect 27246 30036 27252 30048
rect 26660 30008 27252 30036
rect 26660 29996 26666 30008
rect 27246 29996 27252 30008
rect 27304 30036 27310 30048
rect 27430 30036 27436 30048
rect 27304 30008 27436 30036
rect 27304 29996 27310 30008
rect 27430 29996 27436 30008
rect 27488 29996 27494 30048
rect 27522 29996 27528 30048
rect 27580 30036 27586 30048
rect 28721 30039 28779 30045
rect 28721 30036 28733 30039
rect 27580 30008 28733 30036
rect 27580 29996 27586 30008
rect 28721 30005 28733 30008
rect 28767 30005 28779 30039
rect 29104 30036 29132 30203
rect 37550 30200 37556 30212
rect 37608 30200 37614 30252
rect 30098 30172 30104 30184
rect 30059 30144 30104 30172
rect 30098 30132 30104 30144
rect 30156 30132 30162 30184
rect 33321 30175 33379 30181
rect 33321 30141 33333 30175
rect 33367 30141 33379 30175
rect 34238 30172 34244 30184
rect 34199 30144 34244 30172
rect 33321 30135 33379 30141
rect 29270 30104 29276 30116
rect 29231 30076 29276 30104
rect 29270 30064 29276 30076
rect 29328 30064 29334 30116
rect 31573 30107 31631 30113
rect 31573 30073 31585 30107
rect 31619 30104 31631 30107
rect 31662 30104 31668 30116
rect 31619 30076 31668 30104
rect 31619 30073 31631 30076
rect 31573 30067 31631 30073
rect 31662 30064 31668 30076
rect 31720 30064 31726 30116
rect 32398 30104 32404 30116
rect 32359 30076 32404 30104
rect 32398 30064 32404 30076
rect 32456 30064 32462 30116
rect 32582 30064 32588 30116
rect 32640 30104 32646 30116
rect 33336 30104 33364 30135
rect 34238 30132 34244 30144
rect 34296 30132 34302 30184
rect 34348 30144 36032 30172
rect 33778 30104 33784 30116
rect 32640 30076 33784 30104
rect 32640 30064 32646 30076
rect 33778 30064 33784 30076
rect 33836 30104 33842 30116
rect 34348 30104 34376 30144
rect 36004 30113 36032 30144
rect 33836 30076 34376 30104
rect 35989 30107 36047 30113
rect 33836 30064 33842 30076
rect 35989 30073 36001 30107
rect 36035 30073 36047 30107
rect 35989 30067 36047 30073
rect 31386 30036 31392 30048
rect 29104 30008 31392 30036
rect 28721 29999 28779 30005
rect 31386 29996 31392 30008
rect 31444 29996 31450 30048
rect 31754 29996 31760 30048
rect 31812 30036 31818 30048
rect 32600 30036 32628 30064
rect 31812 30008 32628 30036
rect 33413 30039 33471 30045
rect 31812 29996 31818 30008
rect 33413 30005 33425 30039
rect 33459 30036 33471 30039
rect 34606 30036 34612 30048
rect 33459 30008 34612 30036
rect 33459 30005 33471 30008
rect 33413 29999 33471 30005
rect 34606 29996 34612 30008
rect 34664 29996 34670 30048
rect 36538 30036 36544 30048
rect 36499 30008 36544 30036
rect 36538 29996 36544 30008
rect 36596 29996 36602 30048
rect 37458 30036 37464 30048
rect 37419 30008 37464 30036
rect 37458 29996 37464 30008
rect 37516 29996 37522 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 4433 29835 4491 29841
rect 4433 29801 4445 29835
rect 4479 29832 4491 29835
rect 4890 29832 4896 29844
rect 4479 29804 4896 29832
rect 4479 29801 4491 29804
rect 4433 29795 4491 29801
rect 4890 29792 4896 29804
rect 4948 29792 4954 29844
rect 12802 29832 12808 29844
rect 11532 29804 12808 29832
rect 7466 29696 7472 29708
rect 7300 29668 7472 29696
rect 4798 29588 4804 29640
rect 4856 29588 4862 29640
rect 6178 29588 6184 29640
rect 6236 29628 6242 29640
rect 6236 29600 6281 29628
rect 6236 29588 6242 29600
rect 7006 29588 7012 29640
rect 7064 29628 7070 29640
rect 7300 29637 7328 29668
rect 7466 29656 7472 29668
rect 7524 29656 7530 29708
rect 9122 29656 9128 29708
rect 9180 29696 9186 29708
rect 10689 29699 10747 29705
rect 10689 29696 10701 29699
rect 9180 29668 10701 29696
rect 9180 29656 9186 29668
rect 10689 29665 10701 29668
rect 10735 29696 10747 29699
rect 11054 29696 11060 29708
rect 10735 29668 11060 29696
rect 10735 29665 10747 29668
rect 10689 29659 10747 29665
rect 11054 29656 11060 29668
rect 11112 29656 11118 29708
rect 7193 29631 7251 29637
rect 7193 29628 7205 29631
rect 7064 29600 7205 29628
rect 7064 29588 7070 29600
rect 7193 29597 7205 29600
rect 7239 29597 7251 29631
rect 7193 29591 7251 29597
rect 7285 29631 7343 29637
rect 7285 29597 7297 29631
rect 7331 29597 7343 29631
rect 7558 29628 7564 29640
rect 7519 29600 7564 29628
rect 7285 29591 7343 29597
rect 7558 29588 7564 29600
rect 7616 29588 7622 29640
rect 11330 29628 11336 29640
rect 11291 29600 11336 29628
rect 11330 29588 11336 29600
rect 11388 29588 11394 29640
rect 11532 29637 11560 29804
rect 12802 29792 12808 29804
rect 12860 29792 12866 29844
rect 12897 29835 12955 29841
rect 12897 29801 12909 29835
rect 12943 29832 12955 29835
rect 13446 29832 13452 29844
rect 12943 29804 13452 29832
rect 12943 29801 12955 29804
rect 12897 29795 12955 29801
rect 13446 29792 13452 29804
rect 13504 29792 13510 29844
rect 14737 29835 14795 29841
rect 14737 29801 14749 29835
rect 14783 29832 14795 29835
rect 15746 29832 15752 29844
rect 14783 29804 15752 29832
rect 14783 29801 14795 29804
rect 14737 29795 14795 29801
rect 15746 29792 15752 29804
rect 15804 29792 15810 29844
rect 23109 29835 23167 29841
rect 23109 29801 23121 29835
rect 23155 29832 23167 29835
rect 24854 29832 24860 29844
rect 23155 29804 24860 29832
rect 23155 29801 23167 29804
rect 23109 29795 23167 29801
rect 24854 29792 24860 29804
rect 24912 29792 24918 29844
rect 25406 29792 25412 29844
rect 25464 29832 25470 29844
rect 25501 29835 25559 29841
rect 25501 29832 25513 29835
rect 25464 29804 25513 29832
rect 25464 29792 25470 29804
rect 25501 29801 25513 29804
rect 25547 29801 25559 29835
rect 26786 29832 26792 29844
rect 26747 29804 26792 29832
rect 25501 29795 25559 29801
rect 26786 29792 26792 29804
rect 26844 29792 26850 29844
rect 26970 29832 26976 29844
rect 26931 29804 26976 29832
rect 26970 29792 26976 29804
rect 27028 29792 27034 29844
rect 27982 29832 27988 29844
rect 27181 29804 27844 29832
rect 27943 29804 27988 29832
rect 12342 29764 12348 29776
rect 12303 29736 12348 29764
rect 12342 29724 12348 29736
rect 12400 29724 12406 29776
rect 12618 29764 12624 29776
rect 12452 29736 12624 29764
rect 12452 29696 12480 29736
rect 12618 29724 12624 29736
rect 12676 29764 12682 29776
rect 13357 29767 13415 29773
rect 13357 29764 13369 29767
rect 12676 29736 13369 29764
rect 12676 29724 12682 29736
rect 13357 29733 13369 29736
rect 13403 29733 13415 29767
rect 13357 29727 13415 29733
rect 13630 29724 13636 29776
rect 13688 29764 13694 29776
rect 14921 29767 14979 29773
rect 13688 29736 14872 29764
rect 13688 29724 13694 29736
rect 11808 29668 12480 29696
rect 11808 29637 11836 29668
rect 13446 29656 13452 29708
rect 13504 29696 13510 29708
rect 14553 29699 14611 29705
rect 14553 29696 14565 29699
rect 13504 29668 14565 29696
rect 13504 29656 13510 29668
rect 14553 29665 14565 29668
rect 14599 29665 14611 29699
rect 14844 29696 14872 29736
rect 14921 29733 14933 29767
rect 14967 29764 14979 29767
rect 18233 29767 18291 29773
rect 18233 29764 18245 29767
rect 14967 29736 18245 29764
rect 14967 29733 14979 29736
rect 14921 29727 14979 29733
rect 18233 29733 18245 29736
rect 18279 29733 18291 29767
rect 26804 29764 26832 29792
rect 27181 29764 27209 29804
rect 27706 29764 27712 29776
rect 26804 29736 27209 29764
rect 27264 29736 27712 29764
rect 18233 29727 18291 29733
rect 15102 29696 15108 29708
rect 14844 29668 15108 29696
rect 14553 29659 14611 29665
rect 15102 29656 15108 29668
rect 15160 29696 15166 29708
rect 15933 29699 15991 29705
rect 15933 29696 15945 29699
rect 15160 29668 15945 29696
rect 15160 29656 15166 29668
rect 15933 29665 15945 29668
rect 15979 29665 15991 29699
rect 18322 29696 18328 29708
rect 18283 29668 18328 29696
rect 15933 29659 15991 29665
rect 18322 29656 18328 29668
rect 18380 29656 18386 29708
rect 20162 29696 20168 29708
rect 18432 29668 20168 29696
rect 11517 29631 11575 29637
rect 11517 29597 11529 29631
rect 11563 29597 11575 29631
rect 11517 29591 11575 29597
rect 11793 29631 11851 29637
rect 11793 29597 11805 29631
rect 11839 29597 11851 29631
rect 12529 29631 12587 29637
rect 12529 29628 12541 29631
rect 11793 29591 11851 29597
rect 12452 29600 12541 29628
rect 5905 29563 5963 29569
rect 5905 29529 5917 29563
rect 5951 29560 5963 29563
rect 7377 29563 7435 29569
rect 5951 29532 7052 29560
rect 5951 29529 5963 29532
rect 5905 29523 5963 29529
rect 7024 29501 7052 29532
rect 7377 29529 7389 29563
rect 7423 29560 7435 29563
rect 8018 29560 8024 29572
rect 7423 29532 8024 29560
rect 7423 29529 7435 29532
rect 7377 29523 7435 29529
rect 8018 29520 8024 29532
rect 8076 29520 8082 29572
rect 8570 29520 8576 29572
rect 8628 29560 8634 29572
rect 10413 29563 10471 29569
rect 8628 29532 9246 29560
rect 8628 29520 8634 29532
rect 10413 29529 10425 29563
rect 10459 29560 10471 29563
rect 11149 29563 11207 29569
rect 11149 29560 11161 29563
rect 10459 29532 11161 29560
rect 10459 29529 10471 29532
rect 10413 29523 10471 29529
rect 11149 29529 11161 29532
rect 11195 29529 11207 29563
rect 11422 29560 11428 29572
rect 11383 29532 11428 29560
rect 11149 29523 11207 29529
rect 11422 29520 11428 29532
rect 11480 29520 11486 29572
rect 11655 29563 11713 29569
rect 11655 29529 11667 29563
rect 11701 29560 11713 29563
rect 12066 29560 12072 29572
rect 11701 29532 12072 29560
rect 11701 29529 11713 29532
rect 11655 29523 11713 29529
rect 12066 29520 12072 29532
rect 12124 29520 12130 29572
rect 12250 29520 12256 29572
rect 12308 29560 12314 29572
rect 12452 29560 12480 29600
rect 12529 29597 12541 29600
rect 12575 29597 12587 29631
rect 12529 29591 12587 29597
rect 12618 29588 12624 29640
rect 12676 29628 12682 29640
rect 12676 29600 12721 29628
rect 12676 29588 12682 29600
rect 12986 29588 12992 29640
rect 13044 29628 13050 29640
rect 13541 29631 13599 29637
rect 13541 29628 13553 29631
rect 13044 29600 13553 29628
rect 13044 29588 13050 29600
rect 13541 29597 13553 29600
rect 13587 29597 13599 29631
rect 13541 29591 13599 29597
rect 13630 29588 13636 29640
rect 13688 29628 13694 29640
rect 14461 29631 14519 29637
rect 14461 29628 14473 29631
rect 13688 29600 14473 29628
rect 13688 29588 13694 29600
rect 14461 29597 14473 29600
rect 14507 29597 14519 29631
rect 14734 29628 14740 29640
rect 14695 29600 14740 29628
rect 14461 29591 14519 29597
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 15010 29588 15016 29640
rect 15068 29628 15074 29640
rect 15654 29628 15660 29640
rect 15068 29600 15660 29628
rect 15068 29588 15074 29600
rect 15654 29588 15660 29600
rect 15712 29588 15718 29640
rect 16209 29631 16267 29637
rect 16209 29597 16221 29631
rect 16255 29628 16267 29631
rect 16390 29628 16396 29640
rect 16255 29600 16396 29628
rect 16255 29597 16267 29600
rect 16209 29591 16267 29597
rect 16390 29588 16396 29600
rect 16448 29588 16454 29640
rect 17218 29588 17224 29640
rect 17276 29628 17282 29640
rect 17405 29631 17463 29637
rect 17405 29628 17417 29631
rect 17276 29600 17417 29628
rect 17276 29588 17282 29600
rect 17405 29597 17417 29600
rect 17451 29597 17463 29631
rect 17954 29628 17960 29640
rect 17915 29600 17960 29628
rect 17405 29591 17463 29597
rect 17954 29588 17960 29600
rect 18012 29588 18018 29640
rect 18138 29637 18144 29640
rect 18104 29631 18144 29637
rect 18104 29597 18116 29631
rect 18104 29591 18144 29597
rect 18138 29588 18144 29591
rect 18196 29588 18202 29640
rect 12308 29532 12480 29560
rect 12308 29520 12314 29532
rect 14182 29520 14188 29572
rect 14240 29560 14246 29572
rect 15028 29560 15056 29588
rect 14240 29532 15056 29560
rect 14240 29520 14246 29532
rect 15378 29520 15384 29572
rect 15436 29560 15442 29572
rect 16114 29560 16120 29572
rect 15436 29532 16120 29560
rect 15436 29520 15442 29532
rect 16114 29520 16120 29532
rect 16172 29520 16178 29572
rect 18432 29560 18460 29668
rect 20162 29656 20168 29668
rect 20220 29656 20226 29708
rect 20806 29696 20812 29708
rect 20767 29668 20812 29696
rect 20806 29656 20812 29668
rect 20864 29656 20870 29708
rect 24394 29656 24400 29708
rect 24452 29696 24458 29708
rect 24452 29668 25820 29696
rect 24452 29656 24458 29668
rect 18690 29588 18696 29640
rect 18748 29628 18754 29640
rect 19245 29631 19303 29637
rect 19245 29628 19257 29631
rect 18748 29600 19257 29628
rect 18748 29588 18754 29600
rect 19245 29597 19257 29600
rect 19291 29597 19303 29631
rect 19245 29591 19303 29597
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 19392 29600 19441 29628
rect 19392 29588 19398 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19610 29628 19616 29640
rect 19571 29600 19616 29628
rect 19429 29591 19487 29597
rect 19610 29588 19616 29600
rect 19668 29588 19674 29640
rect 23017 29631 23075 29637
rect 23017 29597 23029 29631
rect 23063 29628 23075 29631
rect 23382 29628 23388 29640
rect 23063 29600 23388 29628
rect 23063 29597 23075 29600
rect 23017 29591 23075 29597
rect 23382 29588 23388 29600
rect 23440 29588 23446 29640
rect 23658 29628 23664 29640
rect 23619 29600 23664 29628
rect 23658 29588 23664 29600
rect 23716 29588 23722 29640
rect 24949 29631 25007 29637
rect 24949 29597 24961 29631
rect 24995 29628 25007 29631
rect 25406 29628 25412 29640
rect 24995 29600 25412 29628
rect 24995 29597 25007 29600
rect 24949 29591 25007 29597
rect 25406 29588 25412 29600
rect 25464 29588 25470 29640
rect 25516 29637 25544 29668
rect 25501 29631 25559 29637
rect 25501 29597 25513 29631
rect 25547 29597 25559 29631
rect 25501 29591 25559 29597
rect 25685 29631 25743 29637
rect 25685 29597 25697 29631
rect 25731 29597 25743 29631
rect 25792 29628 25820 29668
rect 27264 29628 27292 29736
rect 27706 29724 27712 29736
rect 27764 29724 27770 29776
rect 25792 29600 27292 29628
rect 25685 29591 25743 29597
rect 16224 29532 18460 29560
rect 19521 29563 19579 29569
rect 7009 29495 7067 29501
rect 7009 29461 7021 29495
rect 7055 29461 7067 29495
rect 7009 29455 7067 29461
rect 8941 29495 8999 29501
rect 8941 29461 8953 29495
rect 8987 29492 8999 29495
rect 10226 29492 10232 29504
rect 8987 29464 10232 29492
rect 8987 29461 8999 29464
rect 8941 29455 8999 29461
rect 10226 29452 10232 29464
rect 10284 29492 10290 29504
rect 12434 29492 12440 29504
rect 10284 29464 12440 29492
rect 10284 29452 10290 29464
rect 12434 29452 12440 29464
rect 12492 29452 12498 29504
rect 12713 29495 12771 29501
rect 12713 29461 12725 29495
rect 12759 29492 12771 29495
rect 12894 29492 12900 29504
rect 12759 29464 12900 29492
rect 12759 29461 12771 29464
rect 12713 29455 12771 29461
rect 12894 29452 12900 29464
rect 12952 29452 12958 29504
rect 15930 29452 15936 29504
rect 15988 29492 15994 29504
rect 16224 29492 16252 29532
rect 19521 29529 19533 29563
rect 19567 29529 19579 29563
rect 21082 29560 21088 29572
rect 21043 29532 21088 29560
rect 19521 29523 19579 29529
rect 17310 29492 17316 29504
rect 15988 29464 16252 29492
rect 17271 29464 17316 29492
rect 15988 29452 15994 29464
rect 17310 29452 17316 29464
rect 17368 29452 17374 29504
rect 18601 29495 18659 29501
rect 18601 29461 18613 29495
rect 18647 29492 18659 29495
rect 19150 29492 19156 29504
rect 18647 29464 19156 29492
rect 18647 29461 18659 29464
rect 18601 29455 18659 29461
rect 19150 29452 19156 29464
rect 19208 29452 19214 29504
rect 19242 29452 19248 29504
rect 19300 29492 19306 29504
rect 19536 29492 19564 29523
rect 21082 29520 21088 29532
rect 21140 29520 21146 29572
rect 22646 29560 22652 29572
rect 22310 29532 22652 29560
rect 22646 29520 22652 29532
rect 22704 29520 22710 29572
rect 25700 29560 25728 29591
rect 27338 29588 27344 29640
rect 27396 29628 27402 29640
rect 27433 29631 27491 29637
rect 27433 29628 27445 29631
rect 27396 29600 27445 29628
rect 27396 29588 27402 29600
rect 27433 29597 27445 29600
rect 27479 29597 27491 29631
rect 27614 29628 27620 29640
rect 27575 29600 27620 29628
rect 27433 29591 27491 29597
rect 27614 29588 27620 29600
rect 27672 29588 27678 29640
rect 27816 29637 27844 29804
rect 27982 29792 27988 29804
rect 28040 29792 28046 29844
rect 28258 29792 28264 29844
rect 28316 29832 28322 29844
rect 28445 29835 28503 29841
rect 28445 29832 28457 29835
rect 28316 29804 28457 29832
rect 28316 29792 28322 29804
rect 28445 29801 28457 29804
rect 28491 29801 28503 29835
rect 28445 29795 28503 29801
rect 28629 29835 28687 29841
rect 28629 29801 28641 29835
rect 28675 29832 28687 29835
rect 28902 29832 28908 29844
rect 28675 29804 28908 29832
rect 28675 29801 28687 29804
rect 28629 29795 28687 29801
rect 28166 29724 28172 29776
rect 28224 29764 28230 29776
rect 28644 29764 28672 29795
rect 28902 29792 28908 29804
rect 28960 29832 28966 29844
rect 29270 29832 29276 29844
rect 28960 29804 29276 29832
rect 28960 29792 28966 29804
rect 29270 29792 29276 29804
rect 29328 29792 29334 29844
rect 30098 29832 30104 29844
rect 30059 29804 30104 29832
rect 30098 29792 30104 29804
rect 30156 29792 30162 29844
rect 32030 29832 32036 29844
rect 31404 29804 32036 29832
rect 28224 29736 28672 29764
rect 28224 29724 28230 29736
rect 29914 29724 29920 29776
rect 29972 29764 29978 29776
rect 30282 29764 30288 29776
rect 29972 29736 30288 29764
rect 29972 29724 29978 29736
rect 30282 29724 30288 29736
rect 30340 29724 30346 29776
rect 31018 29764 31024 29776
rect 30392 29736 31024 29764
rect 30392 29637 30420 29736
rect 31018 29724 31024 29736
rect 31076 29724 31082 29776
rect 31297 29699 31355 29705
rect 31297 29696 31309 29699
rect 30484 29668 31309 29696
rect 30484 29637 30512 29668
rect 31297 29665 31309 29668
rect 31343 29696 31355 29699
rect 31404 29696 31432 29804
rect 32030 29792 32036 29804
rect 32088 29832 32094 29844
rect 32585 29835 32643 29841
rect 32585 29832 32597 29835
rect 32088 29804 32597 29832
rect 32088 29792 32094 29804
rect 32585 29801 32597 29804
rect 32631 29832 32643 29835
rect 32950 29832 32956 29844
rect 32631 29804 32956 29832
rect 32631 29801 32643 29804
rect 32585 29795 32643 29801
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 33502 29792 33508 29844
rect 33560 29832 33566 29844
rect 33873 29835 33931 29841
rect 33873 29832 33885 29835
rect 33560 29804 33885 29832
rect 33560 29792 33566 29804
rect 33873 29801 33885 29804
rect 33919 29801 33931 29835
rect 33873 29795 33931 29801
rect 31941 29767 31999 29773
rect 31941 29733 31953 29767
rect 31987 29733 31999 29767
rect 31941 29727 31999 29733
rect 31343 29668 31432 29696
rect 31343 29665 31355 29668
rect 31297 29659 31355 29665
rect 31478 29656 31484 29708
rect 31536 29696 31542 29708
rect 31956 29696 31984 29727
rect 31536 29668 31581 29696
rect 31956 29668 34100 29696
rect 31536 29656 31542 29668
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29597 27859 29631
rect 27801 29591 27859 29597
rect 30285 29631 30343 29637
rect 30285 29597 30297 29631
rect 30331 29597 30343 29631
rect 30285 29591 30343 29597
rect 30377 29631 30435 29637
rect 30377 29597 30389 29631
rect 30423 29597 30435 29631
rect 30377 29591 30435 29597
rect 30469 29631 30527 29637
rect 30469 29597 30481 29631
rect 30515 29597 30527 29631
rect 30469 29591 30527 29597
rect 30745 29631 30803 29637
rect 30745 29597 30757 29631
rect 30791 29628 30803 29631
rect 31662 29628 31668 29640
rect 30791 29600 31668 29628
rect 30791 29597 30803 29600
rect 30745 29591 30803 29597
rect 26050 29560 26056 29572
rect 25700 29532 26056 29560
rect 26050 29520 26056 29532
rect 26108 29520 26114 29572
rect 26602 29560 26608 29572
rect 26563 29532 26608 29560
rect 26602 29520 26608 29532
rect 26660 29520 26666 29572
rect 26821 29563 26879 29569
rect 26821 29529 26833 29563
rect 26867 29560 26879 29563
rect 27522 29560 27528 29572
rect 26867 29532 27528 29560
rect 26867 29529 26879 29532
rect 26821 29523 26879 29529
rect 27522 29520 27528 29532
rect 27580 29520 27586 29572
rect 27709 29563 27767 29569
rect 27709 29529 27721 29563
rect 27755 29560 27767 29563
rect 27890 29560 27896 29572
rect 27755 29532 27896 29560
rect 27755 29529 27767 29532
rect 27709 29523 27767 29529
rect 27890 29520 27896 29532
rect 27948 29520 27954 29572
rect 28810 29560 28816 29572
rect 28771 29532 28816 29560
rect 28810 29520 28816 29532
rect 28868 29520 28874 29572
rect 19300 29464 19564 29492
rect 19797 29495 19855 29501
rect 19300 29452 19306 29464
rect 19797 29461 19809 29495
rect 19843 29492 19855 29495
rect 20990 29492 20996 29504
rect 19843 29464 20996 29492
rect 19843 29461 19855 29464
rect 19797 29455 19855 29461
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 21818 29452 21824 29504
rect 21876 29492 21882 29504
rect 22557 29495 22615 29501
rect 22557 29492 22569 29495
rect 21876 29464 22569 29492
rect 21876 29452 21882 29464
rect 22557 29461 22569 29464
rect 22603 29461 22615 29495
rect 22557 29455 22615 29461
rect 23845 29495 23903 29501
rect 23845 29461 23857 29495
rect 23891 29492 23903 29495
rect 24762 29492 24768 29504
rect 23891 29464 24768 29492
rect 23891 29461 23903 29464
rect 23845 29455 23903 29461
rect 24762 29452 24768 29464
rect 24820 29452 24826 29504
rect 24857 29495 24915 29501
rect 24857 29461 24869 29495
rect 24903 29492 24915 29495
rect 26694 29492 26700 29504
rect 24903 29464 26700 29492
rect 24903 29461 24915 29464
rect 24857 29455 24915 29461
rect 26694 29452 26700 29464
rect 26752 29492 26758 29504
rect 27982 29492 27988 29504
rect 26752 29464 27988 29492
rect 26752 29452 26758 29464
rect 27982 29452 27988 29464
rect 28040 29452 28046 29504
rect 28613 29495 28671 29501
rect 28613 29461 28625 29495
rect 28659 29492 28671 29495
rect 29086 29492 29092 29504
rect 28659 29464 29092 29492
rect 28659 29461 28671 29464
rect 28613 29455 28671 29461
rect 29086 29452 29092 29464
rect 29144 29452 29150 29504
rect 30300 29492 30328 29591
rect 31662 29588 31668 29600
rect 31720 29628 31726 29640
rect 33226 29628 33232 29640
rect 31720 29600 32812 29628
rect 33187 29600 33232 29628
rect 31720 29588 31726 29600
rect 30650 29569 30656 29572
rect 30607 29563 30656 29569
rect 30607 29529 30619 29563
rect 30653 29529 30656 29563
rect 30607 29523 30656 29529
rect 30650 29520 30656 29523
rect 30708 29520 30714 29572
rect 32784 29569 32812 29600
rect 33226 29588 33232 29600
rect 33284 29588 33290 29640
rect 33410 29628 33416 29640
rect 33371 29600 33416 29628
rect 33410 29588 33416 29600
rect 33468 29588 33474 29640
rect 34072 29637 34100 29668
rect 36078 29656 36084 29708
rect 36136 29696 36142 29708
rect 36265 29699 36323 29705
rect 36265 29696 36277 29699
rect 36136 29668 36277 29696
rect 36136 29656 36142 29668
rect 36265 29665 36277 29668
rect 36311 29665 36323 29699
rect 36265 29659 36323 29665
rect 36449 29699 36507 29705
rect 36449 29665 36461 29699
rect 36495 29696 36507 29699
rect 37458 29696 37464 29708
rect 36495 29668 37464 29696
rect 36495 29665 36507 29668
rect 36449 29659 36507 29665
rect 37458 29656 37464 29668
rect 37516 29656 37522 29708
rect 38102 29696 38108 29708
rect 38063 29668 38108 29696
rect 38102 29656 38108 29668
rect 38160 29656 38166 29708
rect 34057 29631 34115 29637
rect 34057 29597 34069 29631
rect 34103 29597 34115 29631
rect 35526 29628 35532 29640
rect 35487 29600 35532 29628
rect 34057 29591 34115 29597
rect 35526 29588 35532 29600
rect 35584 29588 35590 29640
rect 31573 29563 31631 29569
rect 31573 29560 31585 29563
rect 31220 29532 31585 29560
rect 31220 29492 31248 29532
rect 31573 29529 31585 29532
rect 31619 29560 31631 29563
rect 32769 29563 32827 29569
rect 31619 29532 32720 29560
rect 31619 29529 31631 29532
rect 31573 29523 31631 29529
rect 30300 29464 31248 29492
rect 31386 29452 31392 29504
rect 31444 29492 31450 29504
rect 32122 29492 32128 29504
rect 31444 29464 32128 29492
rect 31444 29452 31450 29464
rect 32122 29452 32128 29464
rect 32180 29452 32186 29504
rect 32306 29452 32312 29504
rect 32364 29492 32370 29504
rect 32582 29501 32588 29504
rect 32401 29495 32459 29501
rect 32401 29492 32413 29495
rect 32364 29464 32413 29492
rect 32364 29452 32370 29464
rect 32401 29461 32413 29464
rect 32447 29461 32459 29495
rect 32401 29455 32459 29461
rect 32569 29495 32588 29501
rect 32569 29461 32581 29495
rect 32569 29455 32588 29461
rect 32582 29452 32588 29455
rect 32640 29452 32646 29504
rect 32692 29492 32720 29532
rect 32769 29529 32781 29563
rect 32815 29529 32827 29563
rect 34698 29560 34704 29572
rect 34659 29532 34704 29560
rect 32769 29523 32827 29529
rect 34698 29520 34704 29532
rect 34756 29520 34762 29572
rect 34885 29563 34943 29569
rect 34885 29529 34897 29563
rect 34931 29560 34943 29563
rect 35342 29560 35348 29572
rect 34931 29532 35348 29560
rect 34931 29529 34943 29532
rect 34885 29523 34943 29529
rect 35342 29520 35348 29532
rect 35400 29520 35406 29572
rect 33321 29495 33379 29501
rect 33321 29492 33333 29495
rect 32692 29464 33333 29492
rect 33321 29461 33333 29464
rect 33367 29461 33379 29495
rect 33321 29455 33379 29461
rect 34514 29452 34520 29504
rect 34572 29492 34578 29504
rect 35069 29495 35127 29501
rect 35069 29492 35081 29495
rect 34572 29464 35081 29492
rect 34572 29452 34578 29464
rect 35069 29461 35081 29464
rect 35115 29461 35127 29495
rect 35069 29455 35127 29461
rect 35621 29495 35679 29501
rect 35621 29461 35633 29495
rect 35667 29492 35679 29495
rect 35894 29492 35900 29504
rect 35667 29464 35900 29492
rect 35667 29461 35679 29464
rect 35621 29455 35679 29461
rect 35894 29452 35900 29464
rect 35952 29452 35958 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 7587 29291 7645 29297
rect 7587 29288 7599 29291
rect 6564 29260 7599 29288
rect 6564 29220 6592 29260
rect 7587 29257 7599 29260
rect 7633 29288 7645 29291
rect 7834 29288 7840 29300
rect 7633 29260 7840 29288
rect 7633 29257 7645 29260
rect 7587 29251 7645 29257
rect 7834 29248 7840 29260
rect 7892 29248 7898 29300
rect 8570 29288 8576 29300
rect 8531 29260 8576 29288
rect 8570 29248 8576 29260
rect 8628 29248 8634 29300
rect 10873 29291 10931 29297
rect 10873 29257 10885 29291
rect 10919 29288 10931 29291
rect 11514 29288 11520 29300
rect 10919 29260 11520 29288
rect 10919 29257 10931 29260
rect 10873 29251 10931 29257
rect 11514 29248 11520 29260
rect 11572 29288 11578 29300
rect 12250 29288 12256 29300
rect 11572 29260 12256 29288
rect 11572 29248 11578 29260
rect 12250 29248 12256 29260
rect 12308 29288 12314 29300
rect 12894 29288 12900 29300
rect 12308 29260 12900 29288
rect 12308 29248 12314 29260
rect 12894 29248 12900 29260
rect 12952 29248 12958 29300
rect 15562 29288 15568 29300
rect 14476 29260 15568 29288
rect 7374 29220 7380 29232
rect 6472 29192 6592 29220
rect 7335 29192 7380 29220
rect 6472 29093 6500 29192
rect 7374 29180 7380 29192
rect 7432 29180 7438 29232
rect 10134 29180 10140 29232
rect 10192 29180 10198 29232
rect 11054 29180 11060 29232
rect 11112 29220 11118 29232
rect 12621 29223 12679 29229
rect 12621 29220 12633 29223
rect 11112 29192 12633 29220
rect 11112 29180 11118 29192
rect 12621 29189 12633 29192
rect 12667 29189 12679 29223
rect 12621 29183 12679 29189
rect 12805 29223 12863 29229
rect 12805 29189 12817 29223
rect 12851 29220 12863 29223
rect 14366 29220 14372 29232
rect 12851 29192 14372 29220
rect 12851 29189 12863 29192
rect 12805 29183 12863 29189
rect 14366 29180 14372 29192
rect 14424 29180 14430 29232
rect 14476 29229 14504 29260
rect 15562 29248 15568 29260
rect 15620 29248 15626 29300
rect 15746 29248 15752 29300
rect 15804 29288 15810 29300
rect 15933 29291 15991 29297
rect 15933 29288 15945 29291
rect 15804 29260 15945 29288
rect 15804 29248 15810 29260
rect 15933 29257 15945 29260
rect 15979 29257 15991 29291
rect 18046 29288 18052 29300
rect 18007 29260 18052 29288
rect 15933 29251 15991 29257
rect 18046 29248 18052 29260
rect 18104 29248 18110 29300
rect 18417 29291 18475 29297
rect 18417 29257 18429 29291
rect 18463 29288 18475 29291
rect 18598 29288 18604 29300
rect 18463 29260 18604 29288
rect 18463 29257 18475 29260
rect 18417 29251 18475 29257
rect 18598 29248 18604 29260
rect 18656 29288 18662 29300
rect 19058 29288 19064 29300
rect 18656 29260 19064 29288
rect 18656 29248 18662 29260
rect 19058 29248 19064 29260
rect 19116 29248 19122 29300
rect 20809 29291 20867 29297
rect 20809 29257 20821 29291
rect 20855 29288 20867 29291
rect 21082 29288 21088 29300
rect 20855 29260 21088 29288
rect 20855 29257 20867 29260
rect 20809 29251 20867 29257
rect 21082 29248 21088 29260
rect 21140 29248 21146 29300
rect 23474 29248 23480 29300
rect 23532 29288 23538 29300
rect 24305 29291 24363 29297
rect 24305 29288 24317 29291
rect 23532 29260 24317 29288
rect 23532 29248 23538 29260
rect 24305 29257 24317 29260
rect 24351 29257 24363 29291
rect 24305 29251 24363 29257
rect 24762 29248 24768 29300
rect 24820 29288 24826 29300
rect 26329 29291 26387 29297
rect 26329 29288 26341 29291
rect 24820 29260 26341 29288
rect 24820 29248 24826 29260
rect 26329 29257 26341 29260
rect 26375 29288 26387 29291
rect 26375 29260 27108 29288
rect 26375 29257 26387 29260
rect 26329 29251 26387 29257
rect 14461 29223 14519 29229
rect 14461 29189 14473 29223
rect 14507 29189 14519 29223
rect 14461 29183 14519 29189
rect 14553 29223 14611 29229
rect 14553 29189 14565 29223
rect 14599 29220 14611 29223
rect 14734 29220 14740 29232
rect 14599 29192 14740 29220
rect 14599 29189 14611 29192
rect 14553 29183 14611 29189
rect 14734 29180 14740 29192
rect 14792 29220 14798 29232
rect 15286 29220 15292 29232
rect 14792 29192 15292 29220
rect 14792 29180 14798 29192
rect 15286 29180 15292 29192
rect 15344 29220 15350 29232
rect 15838 29220 15844 29232
rect 15344 29192 15844 29220
rect 15344 29180 15350 29192
rect 15838 29180 15844 29192
rect 15896 29180 15902 29232
rect 16022 29180 16028 29232
rect 16080 29220 16086 29232
rect 16080 29192 19196 29220
rect 16080 29180 16086 29192
rect 6549 29155 6607 29161
rect 6549 29121 6561 29155
rect 6595 29152 6607 29155
rect 7466 29152 7472 29164
rect 6595 29124 7472 29152
rect 6595 29121 6607 29124
rect 6549 29115 6607 29121
rect 7466 29112 7472 29124
rect 7524 29112 7530 29164
rect 8478 29152 8484 29164
rect 8439 29124 8484 29152
rect 8478 29112 8484 29124
rect 8536 29112 8542 29164
rect 11238 29112 11244 29164
rect 11296 29152 11302 29164
rect 11790 29152 11796 29164
rect 11296 29124 11652 29152
rect 11751 29124 11796 29152
rect 11296 29112 11302 29124
rect 6457 29087 6515 29093
rect 6457 29053 6469 29087
rect 6503 29053 6515 29087
rect 6457 29047 6515 29053
rect 6917 29087 6975 29093
rect 6917 29053 6929 29087
rect 6963 29084 6975 29087
rect 7558 29084 7564 29096
rect 6963 29056 7564 29084
rect 6963 29053 6975 29056
rect 6917 29047 6975 29053
rect 7558 29044 7564 29056
rect 7616 29044 7622 29096
rect 9122 29084 9128 29096
rect 9035 29056 9128 29084
rect 9122 29044 9128 29056
rect 9180 29044 9186 29096
rect 9401 29087 9459 29093
rect 9401 29053 9413 29087
rect 9447 29084 9459 29087
rect 9447 29056 11560 29084
rect 9447 29053 9459 29056
rect 9401 29047 9459 29053
rect 6178 28976 6184 29028
rect 6236 29016 6242 29028
rect 9140 29016 9168 29044
rect 11532 29025 11560 29056
rect 6236 28988 9168 29016
rect 11517 29019 11575 29025
rect 6236 28976 6242 28988
rect 11517 28985 11529 29019
rect 11563 28985 11575 29019
rect 11624 29016 11652 29124
rect 11790 29112 11796 29124
rect 11848 29112 11854 29164
rect 12161 29155 12219 29161
rect 12161 29121 12173 29155
rect 12207 29152 12219 29155
rect 12250 29152 12256 29164
rect 12207 29124 12256 29152
rect 12207 29121 12219 29124
rect 12161 29115 12219 29121
rect 12250 29112 12256 29124
rect 12308 29112 12314 29164
rect 12434 29112 12440 29164
rect 12492 29152 12498 29164
rect 12986 29152 12992 29164
rect 12492 29124 12992 29152
rect 12492 29112 12498 29124
rect 12986 29112 12992 29124
rect 13044 29112 13050 29164
rect 13633 29155 13691 29161
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13814 29152 13820 29164
rect 13775 29124 13820 29152
rect 13633 29115 13691 29121
rect 11701 29087 11759 29093
rect 11701 29053 11713 29087
rect 11747 29084 11759 29087
rect 11974 29084 11980 29096
rect 11747 29056 11980 29084
rect 11747 29053 11759 29056
rect 11701 29047 11759 29053
rect 11974 29044 11980 29056
rect 12032 29044 12038 29096
rect 12069 29087 12127 29093
rect 12069 29053 12081 29087
rect 12115 29053 12127 29087
rect 12069 29047 12127 29053
rect 12084 29016 12112 29047
rect 11624 28988 12112 29016
rect 13648 29016 13676 29115
rect 13814 29112 13820 29124
rect 13872 29112 13878 29164
rect 14277 29155 14335 29161
rect 14277 29121 14289 29155
rect 14323 29121 14335 29155
rect 14277 29115 14335 29121
rect 13725 29087 13783 29093
rect 13725 29053 13737 29087
rect 13771 29084 13783 29087
rect 14292 29084 14320 29115
rect 14642 29112 14648 29164
rect 14700 29152 14706 29164
rect 14700 29124 14745 29152
rect 14700 29112 14706 29124
rect 15654 29112 15660 29164
rect 15712 29152 15718 29164
rect 15749 29155 15807 29161
rect 15749 29152 15761 29155
rect 15712 29124 15761 29152
rect 15712 29112 15718 29124
rect 15749 29121 15761 29124
rect 15795 29121 15807 29155
rect 15749 29115 15807 29121
rect 16117 29155 16175 29161
rect 16117 29121 16129 29155
rect 16163 29152 16175 29155
rect 16206 29152 16212 29164
rect 16163 29124 16212 29152
rect 16163 29121 16175 29124
rect 16117 29115 16175 29121
rect 16206 29112 16212 29124
rect 16264 29152 16270 29164
rect 16482 29152 16488 29164
rect 16264 29124 16488 29152
rect 16264 29112 16270 29124
rect 16482 29112 16488 29124
rect 16540 29152 16546 29164
rect 16669 29155 16727 29161
rect 16669 29152 16681 29155
rect 16540 29124 16681 29152
rect 16540 29112 16546 29124
rect 16669 29121 16681 29124
rect 16715 29121 16727 29155
rect 16669 29115 16727 29121
rect 16945 29155 17003 29161
rect 16945 29121 16957 29155
rect 16991 29121 17003 29155
rect 16945 29115 17003 29121
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29152 17371 29155
rect 17402 29152 17408 29164
rect 17359 29124 17408 29152
rect 17359 29121 17371 29124
rect 17313 29115 17371 29121
rect 13771 29056 14320 29084
rect 13771 29053 13783 29056
rect 13725 29047 13783 29053
rect 15102 29044 15108 29096
rect 15160 29084 15166 29096
rect 16960 29084 16988 29115
rect 17402 29112 17408 29124
rect 17460 29152 17466 29164
rect 18233 29155 18291 29161
rect 18233 29152 18245 29155
rect 17460 29124 18245 29152
rect 17460 29112 17466 29124
rect 18233 29121 18245 29124
rect 18279 29121 18291 29155
rect 18233 29115 18291 29121
rect 18322 29112 18328 29164
rect 18380 29152 18386 29164
rect 18380 29124 18425 29152
rect 18380 29112 18386 29124
rect 15160 29056 16988 29084
rect 18340 29084 18368 29112
rect 19061 29087 19119 29093
rect 19061 29084 19073 29087
rect 18340 29056 19073 29084
rect 15160 29044 15166 29056
rect 19061 29053 19073 29056
rect 19107 29053 19119 29087
rect 19168 29084 19196 29192
rect 23566 29180 23572 29232
rect 23624 29220 23630 29232
rect 24213 29223 24271 29229
rect 24213 29220 24225 29223
rect 23624 29192 24225 29220
rect 23624 29180 23630 29192
rect 24213 29189 24225 29192
rect 24259 29220 24271 29223
rect 24670 29220 24676 29232
rect 24259 29192 24676 29220
rect 24259 29189 24271 29192
rect 24213 29183 24271 29189
rect 24670 29180 24676 29192
rect 24728 29220 24734 29232
rect 25038 29220 25044 29232
rect 24728 29192 25044 29220
rect 24728 29180 24734 29192
rect 25038 29180 25044 29192
rect 25096 29180 25102 29232
rect 25498 29220 25504 29232
rect 25459 29192 25504 29220
rect 25498 29180 25504 29192
rect 25556 29180 25562 29232
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 19337 29155 19395 29161
rect 19337 29152 19349 29155
rect 19300 29124 19349 29152
rect 19300 29112 19306 29124
rect 19337 29121 19349 29124
rect 19383 29121 19395 29155
rect 19337 29115 19395 29121
rect 20898 29112 20904 29164
rect 20956 29152 20962 29164
rect 20993 29155 21051 29161
rect 20993 29152 21005 29155
rect 20956 29124 21005 29152
rect 20956 29112 20962 29124
rect 20993 29121 21005 29124
rect 21039 29121 21051 29155
rect 20993 29115 21051 29121
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29152 21327 29155
rect 21818 29152 21824 29164
rect 21315 29124 21824 29152
rect 21315 29121 21327 29124
rect 21269 29115 21327 29121
rect 21818 29112 21824 29124
rect 21876 29112 21882 29164
rect 25590 29112 25596 29164
rect 25648 29152 25654 29164
rect 26050 29152 26056 29164
rect 25648 29124 26056 29152
rect 25648 29112 25654 29124
rect 26050 29112 26056 29124
rect 26108 29152 26114 29164
rect 26145 29155 26203 29161
rect 26145 29152 26157 29155
rect 26108 29124 26157 29152
rect 26108 29112 26114 29124
rect 26145 29121 26157 29124
rect 26191 29121 26203 29155
rect 26145 29115 26203 29121
rect 26421 29155 26479 29161
rect 26421 29121 26433 29155
rect 26467 29152 26479 29155
rect 26970 29152 26976 29164
rect 26467 29124 26976 29152
rect 26467 29121 26479 29124
rect 26421 29115 26479 29121
rect 26970 29112 26976 29124
rect 27028 29112 27034 29164
rect 27080 29152 27108 29260
rect 27154 29248 27160 29300
rect 27212 29288 27218 29300
rect 27341 29291 27399 29297
rect 27341 29288 27353 29291
rect 27212 29260 27353 29288
rect 27212 29248 27218 29260
rect 27341 29257 27353 29260
rect 27387 29257 27399 29291
rect 27341 29251 27399 29257
rect 27706 29248 27712 29300
rect 27764 29288 27770 29300
rect 28353 29291 28411 29297
rect 28353 29288 28365 29291
rect 27764 29260 28365 29288
rect 27764 29248 27770 29260
rect 28353 29257 28365 29260
rect 28399 29257 28411 29291
rect 28353 29251 28411 29257
rect 28442 29248 28448 29300
rect 28500 29288 28506 29300
rect 29914 29288 29920 29300
rect 28500 29260 29920 29288
rect 28500 29248 28506 29260
rect 29914 29248 29920 29260
rect 29972 29248 29978 29300
rect 30929 29291 30987 29297
rect 30929 29288 30941 29291
rect 30208 29260 30941 29288
rect 27246 29220 27252 29232
rect 27207 29192 27252 29220
rect 27246 29180 27252 29192
rect 27304 29180 27310 29232
rect 29178 29220 29184 29232
rect 28736 29192 29184 29220
rect 27154 29152 27160 29164
rect 27067 29124 27160 29152
rect 27154 29112 27160 29124
rect 27212 29112 27218 29164
rect 28534 29152 28540 29164
rect 28495 29124 28540 29152
rect 28534 29112 28540 29124
rect 28592 29112 28598 29164
rect 28736 29161 28764 29192
rect 29178 29180 29184 29192
rect 29236 29180 29242 29232
rect 28721 29155 28779 29161
rect 28721 29121 28733 29155
rect 28767 29121 28779 29155
rect 28721 29115 28779 29121
rect 28810 29112 28816 29164
rect 28868 29152 28874 29164
rect 29089 29155 29147 29161
rect 29089 29152 29101 29155
rect 28868 29124 29101 29152
rect 28868 29112 28874 29124
rect 29089 29121 29101 29124
rect 29135 29121 29147 29155
rect 29089 29115 29147 29121
rect 29641 29155 29699 29161
rect 29641 29121 29653 29155
rect 29687 29152 29699 29155
rect 30208 29152 30236 29260
rect 30929 29257 30941 29260
rect 30975 29257 30987 29291
rect 30929 29251 30987 29257
rect 31018 29248 31024 29300
rect 31076 29288 31082 29300
rect 32125 29291 32183 29297
rect 32125 29288 32137 29291
rect 31076 29260 32137 29288
rect 31076 29248 31082 29260
rect 32125 29257 32137 29260
rect 32171 29257 32183 29291
rect 32125 29251 32183 29257
rect 32214 29248 32220 29300
rect 32272 29288 32278 29300
rect 32272 29260 33916 29288
rect 32272 29248 32278 29260
rect 31481 29223 31539 29229
rect 31481 29220 31493 29223
rect 30668 29192 31493 29220
rect 29687 29124 30236 29152
rect 30377 29155 30435 29161
rect 29687 29121 29699 29124
rect 29641 29115 29699 29121
rect 30377 29121 30389 29155
rect 30423 29152 30435 29155
rect 30668 29152 30696 29192
rect 31481 29189 31493 29192
rect 31527 29220 31539 29223
rect 33226 29220 33232 29232
rect 31527 29192 33232 29220
rect 31527 29189 31539 29192
rect 31481 29183 31539 29189
rect 33226 29180 33232 29192
rect 33284 29180 33290 29232
rect 30423 29124 30512 29152
rect 30423 29121 30435 29124
rect 30377 29115 30435 29121
rect 22002 29084 22008 29096
rect 19168 29056 21312 29084
rect 21963 29056 22008 29084
rect 19061 29047 19119 29053
rect 14918 29016 14924 29028
rect 13648 28988 14924 29016
rect 11517 28979 11575 28985
rect 14918 28976 14924 28988
rect 14976 28976 14982 29028
rect 15565 29019 15623 29025
rect 15565 28985 15577 29019
rect 15611 29016 15623 29019
rect 16114 29016 16120 29028
rect 15611 28988 16120 29016
rect 15611 28985 15623 28988
rect 15565 28979 15623 28985
rect 16114 28976 16120 28988
rect 16172 28976 16178 29028
rect 18506 28976 18512 29028
rect 18564 29016 18570 29028
rect 18601 29019 18659 29025
rect 18601 29016 18613 29019
rect 18564 28988 18613 29016
rect 18564 28976 18570 28988
rect 18601 28985 18613 28988
rect 18647 28985 18659 29019
rect 19076 29016 19104 29047
rect 19518 29016 19524 29028
rect 19076 28988 19524 29016
rect 18601 28979 18659 28985
rect 19518 28976 19524 28988
rect 19576 28976 19582 29028
rect 21174 29016 21180 29028
rect 21135 28988 21180 29016
rect 21174 28976 21180 28988
rect 21232 28976 21238 29028
rect 21284 29016 21312 29056
rect 22002 29044 22008 29056
rect 22060 29044 22066 29096
rect 22281 29087 22339 29093
rect 22281 29053 22293 29087
rect 22327 29053 22339 29087
rect 22281 29047 22339 29053
rect 25685 29087 25743 29093
rect 25685 29053 25697 29087
rect 25731 29084 25743 29087
rect 26510 29084 26516 29096
rect 25731 29056 26516 29084
rect 25731 29053 25743 29056
rect 25685 29047 25743 29053
rect 22296 29016 22324 29047
rect 26510 29044 26516 29056
rect 26568 29084 26574 29096
rect 27614 29084 27620 29096
rect 26568 29056 27620 29084
rect 26568 29044 26574 29056
rect 27614 29044 27620 29056
rect 27672 29044 27678 29096
rect 30285 29087 30343 29093
rect 30285 29084 30297 29087
rect 28736 29056 30297 29084
rect 28736 29028 28764 29056
rect 30285 29053 30297 29056
rect 30331 29053 30343 29087
rect 30285 29047 30343 29053
rect 21284 28988 22324 29016
rect 25130 28976 25136 29028
rect 25188 29016 25194 29028
rect 25958 29016 25964 29028
rect 25188 28988 25964 29016
rect 25188 28976 25194 28988
rect 25958 28976 25964 28988
rect 26016 29016 26022 29028
rect 26973 29019 27031 29025
rect 26973 29016 26985 29019
rect 26016 28988 26985 29016
rect 26016 28976 26022 28988
rect 26973 28985 26985 28988
rect 27019 28985 27031 29019
rect 26973 28979 27031 28985
rect 7466 28908 7472 28960
rect 7524 28948 7530 28960
rect 7561 28951 7619 28957
rect 7561 28948 7573 28951
rect 7524 28920 7573 28948
rect 7524 28908 7530 28920
rect 7561 28917 7573 28920
rect 7607 28917 7619 28951
rect 7742 28948 7748 28960
rect 7703 28920 7748 28948
rect 7561 28911 7619 28917
rect 7742 28908 7748 28920
rect 7800 28908 7806 28960
rect 14366 28908 14372 28960
rect 14424 28948 14430 28960
rect 14829 28951 14887 28957
rect 14829 28948 14841 28951
rect 14424 28920 14841 28948
rect 14424 28908 14430 28920
rect 14829 28917 14841 28920
rect 14875 28917 14887 28951
rect 14829 28911 14887 28917
rect 17221 28951 17279 28957
rect 17221 28917 17233 28951
rect 17267 28948 17279 28951
rect 18414 28948 18420 28960
rect 17267 28920 18420 28948
rect 17267 28917 17279 28920
rect 17221 28911 17279 28917
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 26145 28951 26203 28957
rect 26145 28917 26157 28951
rect 26191 28948 26203 28951
rect 26234 28948 26240 28960
rect 26191 28920 26240 28948
rect 26191 28917 26203 28920
rect 26145 28911 26203 28917
rect 26234 28908 26240 28920
rect 26292 28908 26298 28960
rect 26988 28948 27016 28979
rect 27062 28976 27068 29028
rect 27120 29016 27126 29028
rect 27525 29019 27583 29025
rect 27525 29016 27537 29019
rect 27120 28988 27537 29016
rect 27120 28976 27126 28988
rect 27525 28985 27537 28988
rect 27571 28985 27583 29019
rect 27525 28979 27583 28985
rect 28718 28976 28724 29028
rect 28776 28976 28782 29028
rect 28902 28976 28908 29028
rect 28960 29016 28966 29028
rect 30484 29016 30512 29124
rect 28960 28988 30512 29016
rect 30576 29124 30696 29152
rect 30745 29155 30803 29161
rect 28960 28976 28966 28988
rect 30576 28960 30604 29124
rect 30745 29121 30757 29155
rect 30791 29121 30803 29155
rect 31386 29152 31392 29164
rect 31347 29124 31392 29152
rect 30745 29115 30803 29121
rect 30760 29084 30788 29115
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 31573 29155 31631 29161
rect 31754 29158 31760 29164
rect 31573 29121 31585 29155
rect 31619 29152 31631 29155
rect 31726 29152 31760 29158
rect 31619 29124 31760 29152
rect 31619 29121 31631 29124
rect 31573 29115 31631 29121
rect 31754 29112 31760 29124
rect 31812 29112 31818 29164
rect 32122 29152 32128 29164
rect 32083 29124 32128 29152
rect 32122 29112 32128 29124
rect 32180 29112 32186 29164
rect 32306 29152 32312 29164
rect 32267 29124 32312 29152
rect 32306 29112 32312 29124
rect 32364 29112 32370 29164
rect 32950 29152 32956 29164
rect 32911 29124 32956 29152
rect 32950 29112 32956 29124
rect 33008 29112 33014 29164
rect 33888 29161 33916 29260
rect 36538 29220 36544 29232
rect 36110 29192 36544 29220
rect 36538 29180 36544 29192
rect 36596 29180 36602 29232
rect 33413 29155 33471 29161
rect 33413 29121 33425 29155
rect 33459 29121 33471 29155
rect 33413 29115 33471 29121
rect 33873 29155 33931 29161
rect 33873 29121 33885 29155
rect 33919 29121 33931 29155
rect 33873 29115 33931 29121
rect 32858 29084 32864 29096
rect 30760 29056 32864 29084
rect 32858 29044 32864 29056
rect 32916 29044 32922 29096
rect 33134 29084 33140 29096
rect 33095 29056 33140 29084
rect 33134 29044 33140 29056
rect 33192 29044 33198 29096
rect 33428 29084 33456 29115
rect 34238 29112 34244 29164
rect 34296 29152 34302 29164
rect 34609 29155 34667 29161
rect 34609 29152 34621 29155
rect 34296 29124 34621 29152
rect 34296 29112 34302 29124
rect 34609 29121 34621 29124
rect 34655 29121 34667 29155
rect 37550 29152 37556 29164
rect 37511 29124 37556 29152
rect 34609 29115 34667 29121
rect 37550 29112 37556 29124
rect 37608 29112 37614 29164
rect 33686 29084 33692 29096
rect 33428 29056 33692 29084
rect 33686 29044 33692 29056
rect 33744 29084 33750 29096
rect 35342 29084 35348 29096
rect 33744 29056 35348 29084
rect 33744 29044 33750 29056
rect 35342 29044 35348 29056
rect 35400 29084 35406 29096
rect 36357 29087 36415 29093
rect 36357 29084 36369 29087
rect 35400 29056 36369 29084
rect 35400 29044 35406 29056
rect 36357 29053 36369 29056
rect 36403 29053 36415 29087
rect 36357 29047 36415 29053
rect 32769 29019 32827 29025
rect 32769 29016 32781 29019
rect 30852 28988 32781 29016
rect 27246 28948 27252 28960
rect 26988 28920 27252 28948
rect 27246 28908 27252 28920
rect 27304 28908 27310 28960
rect 30558 28908 30564 28960
rect 30616 28908 30622 28960
rect 30745 28951 30803 28957
rect 30745 28917 30757 28951
rect 30791 28948 30803 28951
rect 30852 28948 30880 28988
rect 32769 28985 32781 28988
rect 32815 28985 32827 29019
rect 32769 28979 32827 28985
rect 30791 28920 30880 28948
rect 30791 28917 30803 28920
rect 30745 28911 30803 28917
rect 30926 28908 30932 28960
rect 30984 28948 30990 28960
rect 31478 28948 31484 28960
rect 30984 28920 31484 28948
rect 30984 28908 30990 28920
rect 31478 28908 31484 28920
rect 31536 28908 31542 28960
rect 33321 28951 33379 28957
rect 33321 28917 33333 28951
rect 33367 28948 33379 28951
rect 33778 28948 33784 28960
rect 33367 28920 33784 28948
rect 33367 28917 33379 28920
rect 33321 28911 33379 28917
rect 33778 28908 33784 28920
rect 33836 28908 33842 28960
rect 33965 28951 34023 28957
rect 33965 28917 33977 28951
rect 34011 28948 34023 28951
rect 34054 28948 34060 28960
rect 34011 28920 34060 28948
rect 34011 28917 34023 28920
rect 33965 28911 34023 28917
rect 34054 28908 34060 28920
rect 34112 28908 34118 28960
rect 34146 28908 34152 28960
rect 34204 28948 34210 28960
rect 34866 28951 34924 28957
rect 34866 28948 34878 28951
rect 34204 28920 34878 28948
rect 34204 28908 34210 28920
rect 34866 28917 34878 28920
rect 34912 28917 34924 28951
rect 34866 28911 34924 28917
rect 37645 28951 37703 28957
rect 37645 28917 37657 28951
rect 37691 28948 37703 28951
rect 37918 28948 37924 28960
rect 37691 28920 37924 28948
rect 37691 28917 37703 28920
rect 37645 28911 37703 28917
rect 37918 28908 37924 28920
rect 37976 28908 37982 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 9125 28747 9183 28753
rect 9125 28713 9137 28747
rect 9171 28744 9183 28747
rect 9950 28744 9956 28756
rect 9171 28716 9956 28744
rect 9171 28713 9183 28716
rect 9125 28707 9183 28713
rect 9950 28704 9956 28716
rect 10008 28704 10014 28756
rect 11330 28704 11336 28756
rect 11388 28744 11394 28756
rect 11701 28747 11759 28753
rect 11701 28744 11713 28747
rect 11388 28716 11713 28744
rect 11388 28704 11394 28716
rect 11701 28713 11713 28716
rect 11747 28713 11759 28747
rect 15838 28744 15844 28756
rect 15799 28716 15844 28744
rect 11701 28707 11759 28713
rect 15838 28704 15844 28716
rect 15896 28704 15902 28756
rect 19518 28744 19524 28756
rect 19479 28716 19524 28744
rect 19518 28704 19524 28716
rect 19576 28704 19582 28756
rect 24397 28747 24455 28753
rect 24397 28713 24409 28747
rect 24443 28744 24455 28747
rect 25130 28744 25136 28756
rect 24443 28716 25136 28744
rect 24443 28713 24455 28716
rect 24397 28707 24455 28713
rect 25130 28704 25136 28716
rect 25188 28704 25194 28756
rect 28718 28704 28724 28756
rect 28776 28744 28782 28756
rect 28813 28747 28871 28753
rect 28813 28744 28825 28747
rect 28776 28716 28825 28744
rect 28776 28704 28782 28716
rect 28813 28713 28825 28716
rect 28859 28713 28871 28747
rect 28994 28744 29000 28756
rect 28955 28716 29000 28744
rect 28813 28707 28871 28713
rect 28994 28704 29000 28716
rect 29052 28704 29058 28756
rect 30466 28744 30472 28756
rect 30427 28716 30472 28744
rect 30466 28704 30472 28716
rect 30524 28704 30530 28756
rect 31018 28744 31024 28756
rect 30944 28716 31024 28744
rect 9769 28679 9827 28685
rect 9769 28645 9781 28679
rect 9815 28676 9827 28679
rect 9858 28676 9864 28688
rect 9815 28648 9864 28676
rect 9815 28645 9827 28648
rect 9769 28639 9827 28645
rect 9858 28636 9864 28648
rect 9916 28676 9922 28688
rect 11146 28676 11152 28688
rect 9916 28648 11152 28676
rect 9916 28636 9922 28648
rect 11146 28636 11152 28648
rect 11204 28636 11210 28688
rect 11422 28636 11428 28688
rect 11480 28676 11486 28688
rect 13081 28679 13139 28685
rect 13081 28676 13093 28679
rect 11480 28648 13093 28676
rect 11480 28636 11486 28648
rect 13081 28645 13093 28648
rect 13127 28645 13139 28679
rect 18690 28676 18696 28688
rect 18651 28648 18696 28676
rect 13081 28639 13139 28645
rect 18690 28636 18696 28648
rect 18748 28636 18754 28688
rect 26878 28636 26884 28688
rect 26936 28636 26942 28688
rect 29822 28676 29828 28688
rect 28644 28648 29828 28676
rect 7374 28608 7380 28620
rect 7335 28580 7380 28608
rect 7374 28568 7380 28580
rect 7432 28568 7438 28620
rect 12618 28608 12624 28620
rect 12406 28580 12624 28608
rect 7098 28540 7104 28552
rect 7059 28512 7104 28540
rect 7098 28500 7104 28512
rect 7156 28500 7162 28552
rect 10226 28500 10232 28552
rect 10284 28540 10290 28552
rect 10781 28543 10839 28549
rect 10781 28540 10793 28543
rect 10284 28512 10793 28540
rect 10284 28500 10290 28512
rect 10781 28509 10793 28512
rect 10827 28509 10839 28543
rect 10781 28503 10839 28509
rect 11885 28543 11943 28549
rect 11885 28509 11897 28543
rect 11931 28540 11943 28543
rect 12406 28540 12434 28580
rect 12618 28568 12624 28580
rect 12676 28608 12682 28620
rect 14093 28611 14151 28617
rect 12676 28580 13216 28608
rect 12676 28568 12682 28580
rect 13188 28549 13216 28580
rect 14093 28577 14105 28611
rect 14139 28608 14151 28611
rect 14458 28608 14464 28620
rect 14139 28580 14464 28608
rect 14139 28577 14151 28580
rect 14093 28571 14151 28577
rect 14458 28568 14464 28580
rect 14516 28568 14522 28620
rect 15378 28568 15384 28620
rect 15436 28608 15442 28620
rect 16393 28611 16451 28617
rect 15436 28580 15608 28608
rect 15436 28568 15442 28580
rect 11931 28512 12434 28540
rect 12989 28543 13047 28549
rect 11931 28509 11943 28512
rect 11885 28503 11943 28509
rect 12989 28509 13001 28543
rect 13035 28509 13047 28543
rect 12989 28503 13047 28509
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28509 13231 28543
rect 15580 28540 15608 28580
rect 16393 28577 16405 28611
rect 16439 28608 16451 28611
rect 17313 28611 17371 28617
rect 17313 28608 17325 28611
rect 16439 28580 17325 28608
rect 16439 28577 16451 28580
rect 16393 28571 16451 28577
rect 17313 28577 17325 28580
rect 17359 28577 17371 28611
rect 17313 28571 17371 28577
rect 17402 28568 17408 28620
rect 17460 28608 17466 28620
rect 17678 28608 17684 28620
rect 17460 28580 17684 28608
rect 17460 28568 17466 28580
rect 17678 28568 17684 28580
rect 17736 28568 17742 28620
rect 18414 28608 18420 28620
rect 18375 28580 18420 28608
rect 18414 28568 18420 28580
rect 18472 28568 18478 28620
rect 20898 28568 20904 28620
rect 20956 28608 20962 28620
rect 21269 28611 21327 28617
rect 21269 28608 21281 28611
rect 20956 28580 21281 28608
rect 20956 28568 20962 28580
rect 21269 28577 21281 28580
rect 21315 28577 21327 28611
rect 23566 28608 23572 28620
rect 23527 28580 23572 28608
rect 21269 28571 21327 28577
rect 23566 28568 23572 28580
rect 23624 28568 23630 28620
rect 26142 28608 26148 28620
rect 26103 28580 26148 28608
rect 26142 28568 26148 28580
rect 26200 28568 26206 28620
rect 26789 28611 26847 28617
rect 26789 28577 26801 28611
rect 26835 28608 26847 28611
rect 26896 28608 26924 28636
rect 26835 28580 28028 28608
rect 26835 28577 26847 28580
rect 26789 28571 26847 28577
rect 16485 28543 16543 28549
rect 16485 28540 16497 28543
rect 15580 28512 16497 28540
rect 13173 28503 13231 28509
rect 16485 28509 16497 28512
rect 16531 28509 16543 28543
rect 16485 28503 16543 28509
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28509 16635 28543
rect 16577 28503 16635 28509
rect 16669 28543 16727 28549
rect 16669 28509 16681 28543
rect 16715 28540 16727 28543
rect 16758 28540 16764 28552
rect 16715 28512 16764 28540
rect 16715 28509 16727 28512
rect 16669 28503 16727 28509
rect 7742 28432 7748 28484
rect 7800 28472 7806 28484
rect 9093 28475 9151 28481
rect 9093 28472 9105 28475
rect 7800 28444 9105 28472
rect 7800 28432 7806 28444
rect 9093 28441 9105 28444
rect 9139 28441 9151 28475
rect 9093 28435 9151 28441
rect 9309 28475 9367 28481
rect 9309 28441 9321 28475
rect 9355 28472 9367 28475
rect 9674 28472 9680 28484
rect 9355 28444 9680 28472
rect 9355 28441 9367 28444
rect 9309 28435 9367 28441
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 9950 28472 9956 28484
rect 9911 28444 9956 28472
rect 9950 28432 9956 28444
rect 10008 28432 10014 28484
rect 8938 28404 8944 28416
rect 8899 28376 8944 28404
rect 8938 28364 8944 28376
rect 8996 28364 9002 28416
rect 10226 28364 10232 28416
rect 10284 28404 10290 28416
rect 10597 28407 10655 28413
rect 10597 28404 10609 28407
rect 10284 28376 10609 28404
rect 10284 28364 10290 28376
rect 10597 28373 10609 28376
rect 10643 28373 10655 28407
rect 10796 28404 10824 28503
rect 11974 28432 11980 28484
rect 12032 28472 12038 28484
rect 12069 28475 12127 28481
rect 12069 28472 12081 28475
rect 12032 28444 12081 28472
rect 12032 28432 12038 28444
rect 12069 28441 12081 28444
rect 12115 28472 12127 28475
rect 13004 28472 13032 28503
rect 14366 28472 14372 28484
rect 12115 28444 13032 28472
rect 14327 28444 14372 28472
rect 12115 28441 12127 28444
rect 12069 28435 12127 28441
rect 14366 28432 14372 28444
rect 14424 28432 14430 28484
rect 15746 28472 15752 28484
rect 15594 28444 15752 28472
rect 15746 28432 15752 28444
rect 15804 28432 15810 28484
rect 16592 28472 16620 28503
rect 16758 28500 16764 28512
rect 16816 28500 16822 28552
rect 17494 28540 17500 28552
rect 17455 28512 17500 28540
rect 17494 28500 17500 28512
rect 17552 28500 17558 28552
rect 18325 28543 18383 28549
rect 18325 28509 18337 28543
rect 18371 28540 18383 28543
rect 18966 28540 18972 28552
rect 18371 28512 18972 28540
rect 18371 28509 18383 28512
rect 18325 28503 18383 28509
rect 18966 28500 18972 28512
rect 19024 28540 19030 28552
rect 19242 28540 19248 28552
rect 19024 28512 19248 28540
rect 19024 28500 19030 28512
rect 19242 28500 19248 28512
rect 19300 28500 19306 28552
rect 21358 28500 21364 28552
rect 21416 28540 21422 28552
rect 21729 28543 21787 28549
rect 21729 28540 21741 28543
rect 21416 28512 21741 28540
rect 21416 28500 21422 28512
rect 21729 28509 21741 28512
rect 21775 28509 21787 28543
rect 22557 28543 22615 28549
rect 22557 28540 22569 28543
rect 21729 28503 21787 28509
rect 22388 28512 22569 28540
rect 18414 28472 18420 28484
rect 16592 28444 18420 28472
rect 18414 28432 18420 28444
rect 18472 28432 18478 28484
rect 20990 28472 20996 28484
rect 20562 28444 20852 28472
rect 20951 28444 20996 28472
rect 12618 28404 12624 28416
rect 10796 28376 12624 28404
rect 10597 28367 10655 28373
rect 12618 28364 12624 28376
rect 12676 28364 12682 28416
rect 12710 28364 12716 28416
rect 12768 28404 12774 28416
rect 16666 28404 16672 28416
rect 12768 28376 16672 28404
rect 12768 28364 12774 28376
rect 16666 28364 16672 28376
rect 16724 28364 16730 28416
rect 16853 28407 16911 28413
rect 16853 28373 16865 28407
rect 16899 28404 16911 28407
rect 16942 28404 16948 28416
rect 16899 28376 16948 28404
rect 16899 28373 16911 28376
rect 16853 28367 16911 28373
rect 16942 28364 16948 28376
rect 17000 28364 17006 28416
rect 20824 28404 20852 28444
rect 20990 28432 20996 28444
rect 21048 28432 21054 28484
rect 21821 28407 21879 28413
rect 21821 28404 21833 28407
rect 20824 28376 21833 28404
rect 21821 28373 21833 28376
rect 21867 28373 21879 28407
rect 22388 28404 22416 28512
rect 22557 28509 22569 28512
rect 22603 28509 22615 28543
rect 22557 28503 22615 28509
rect 22922 28500 22928 28552
rect 22980 28540 22986 28552
rect 23845 28543 23903 28549
rect 23845 28540 23857 28543
rect 22980 28512 23857 28540
rect 22980 28500 22986 28512
rect 23845 28509 23857 28512
rect 23891 28509 23903 28543
rect 26878 28540 26884 28552
rect 26839 28512 26884 28540
rect 23845 28503 23903 28509
rect 26878 28500 26884 28512
rect 26936 28500 26942 28552
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28509 27031 28543
rect 26973 28503 27031 28509
rect 27065 28543 27123 28549
rect 27065 28509 27077 28543
rect 27111 28540 27123 28543
rect 27246 28540 27252 28552
rect 27111 28512 27252 28540
rect 27111 28509 27123 28512
rect 27065 28503 27123 28509
rect 22465 28475 22523 28481
rect 22465 28441 22477 28475
rect 22511 28472 22523 28475
rect 25866 28472 25872 28484
rect 22511 28444 24702 28472
rect 25827 28444 25872 28472
rect 22511 28441 22523 28444
rect 22465 28435 22523 28441
rect 25866 28432 25872 28444
rect 25924 28432 25930 28484
rect 26988 28472 27016 28503
rect 27246 28500 27252 28512
rect 27304 28500 27310 28552
rect 28000 28549 28028 28580
rect 27985 28543 28043 28549
rect 27985 28509 27997 28543
rect 28031 28509 28043 28543
rect 27985 28503 28043 28509
rect 27154 28472 27160 28484
rect 26988 28444 27160 28472
rect 27154 28432 27160 28444
rect 27212 28472 27218 28484
rect 28644 28481 28672 28648
rect 29822 28636 29828 28648
rect 29880 28636 29886 28688
rect 30009 28679 30067 28685
rect 30009 28645 30021 28679
rect 30055 28676 30067 28679
rect 30834 28676 30840 28688
rect 30055 28648 30840 28676
rect 30055 28645 30067 28648
rect 30009 28639 30067 28645
rect 30834 28636 30840 28648
rect 30892 28636 30898 28688
rect 30558 28608 30564 28620
rect 29564 28580 30564 28608
rect 29564 28549 29592 28580
rect 30558 28568 30564 28580
rect 30616 28568 30622 28620
rect 29549 28543 29607 28549
rect 29549 28509 29561 28543
rect 29595 28509 29607 28543
rect 29822 28540 29828 28552
rect 29783 28512 29828 28540
rect 29549 28503 29607 28509
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 30650 28540 30656 28552
rect 30611 28512 30656 28540
rect 30650 28500 30656 28512
rect 30708 28500 30714 28552
rect 30742 28500 30748 28552
rect 30800 28540 30806 28552
rect 30944 28549 30972 28716
rect 31018 28704 31024 28716
rect 31076 28704 31082 28756
rect 31202 28704 31208 28756
rect 31260 28744 31266 28756
rect 31570 28744 31576 28756
rect 31260 28716 31432 28744
rect 31531 28716 31576 28744
rect 31260 28704 31266 28716
rect 31404 28676 31432 28716
rect 31570 28704 31576 28716
rect 31628 28704 31634 28756
rect 31662 28704 31668 28756
rect 31720 28744 31726 28756
rect 33410 28744 33416 28756
rect 31720 28716 33416 28744
rect 31720 28704 31726 28716
rect 33410 28704 33416 28716
rect 33468 28704 33474 28756
rect 34146 28744 34152 28756
rect 34107 28716 34152 28744
rect 34146 28704 34152 28716
rect 34204 28704 34210 28756
rect 34606 28704 34612 28756
rect 34664 28744 34670 28756
rect 35529 28747 35587 28753
rect 35529 28744 35541 28747
rect 34664 28716 35541 28744
rect 34664 28704 34670 28716
rect 35529 28713 35541 28716
rect 35575 28713 35587 28747
rect 35529 28707 35587 28713
rect 31404 28648 31616 28676
rect 31588 28620 31616 28648
rect 33134 28636 33140 28688
rect 33192 28676 33198 28688
rect 33192 28648 35020 28676
rect 33192 28636 33198 28648
rect 31570 28568 31576 28620
rect 31628 28608 31634 28620
rect 31628 28580 33272 28608
rect 31628 28568 31634 28580
rect 30837 28543 30895 28549
rect 30837 28540 30849 28543
rect 30800 28512 30849 28540
rect 30800 28500 30806 28512
rect 30837 28509 30849 28512
rect 30883 28509 30895 28543
rect 30837 28503 30895 28509
rect 30929 28543 30987 28549
rect 30929 28509 30941 28543
rect 30975 28509 30987 28543
rect 30929 28503 30987 28509
rect 31018 28500 31024 28552
rect 31076 28540 31082 28552
rect 31389 28543 31447 28549
rect 31389 28540 31401 28543
rect 31076 28512 31401 28540
rect 31076 28500 31082 28512
rect 31389 28509 31401 28512
rect 31435 28509 31447 28543
rect 32306 28540 32312 28552
rect 31389 28503 31447 28509
rect 31726 28512 32312 28540
rect 27801 28475 27859 28481
rect 27801 28472 27813 28475
rect 27212 28444 27813 28472
rect 27212 28432 27218 28444
rect 27801 28441 27813 28444
rect 27847 28441 27859 28475
rect 27801 28435 27859 28441
rect 28629 28475 28687 28481
rect 28629 28441 28641 28475
rect 28675 28441 28687 28475
rect 28629 28435 28687 28441
rect 28845 28475 28903 28481
rect 28845 28441 28857 28475
rect 28891 28472 28903 28475
rect 31726 28472 31754 28512
rect 32306 28500 32312 28512
rect 32364 28500 32370 28552
rect 33244 28540 33272 28580
rect 33318 28568 33324 28620
rect 33376 28608 33382 28620
rect 33505 28611 33563 28617
rect 33505 28608 33517 28611
rect 33376 28580 33517 28608
rect 33376 28568 33382 28580
rect 33505 28577 33517 28580
rect 33551 28577 33563 28611
rect 34790 28608 34796 28620
rect 33505 28571 33563 28577
rect 33704 28580 34796 28608
rect 33704 28540 33732 28580
rect 34790 28568 34796 28580
rect 34848 28568 34854 28620
rect 34992 28552 35020 28648
rect 35069 28611 35127 28617
rect 35069 28577 35081 28611
rect 35115 28608 35127 28611
rect 35342 28608 35348 28620
rect 35115 28580 35348 28608
rect 35115 28577 35127 28580
rect 35069 28571 35127 28577
rect 35342 28568 35348 28580
rect 35400 28568 35406 28620
rect 37182 28608 37188 28620
rect 37143 28580 37188 28608
rect 37182 28568 37188 28580
rect 37240 28568 37246 28620
rect 37918 28608 37924 28620
rect 37879 28580 37924 28608
rect 37918 28568 37924 28580
rect 37976 28568 37982 28620
rect 33244 28512 33732 28540
rect 33778 28500 33784 28552
rect 33836 28540 33842 28552
rect 33965 28543 34023 28549
rect 33836 28512 33881 28540
rect 33836 28500 33842 28512
rect 33965 28509 33977 28543
rect 34011 28540 34023 28543
rect 34514 28540 34520 28552
rect 34011 28512 34520 28540
rect 34011 28509 34023 28512
rect 33965 28503 34023 28509
rect 34514 28500 34520 28512
rect 34572 28500 34578 28552
rect 34885 28543 34943 28549
rect 34885 28509 34897 28543
rect 34931 28540 34943 28543
rect 34974 28540 34980 28552
rect 34931 28512 34980 28540
rect 34931 28509 34943 28512
rect 34885 28503 34943 28509
rect 34974 28500 34980 28512
rect 35032 28500 35038 28552
rect 35529 28543 35587 28549
rect 35529 28509 35541 28543
rect 35575 28509 35587 28543
rect 35713 28543 35771 28549
rect 35713 28540 35725 28543
rect 35529 28503 35587 28509
rect 35636 28512 35725 28540
rect 28891 28444 31754 28472
rect 32401 28475 32459 28481
rect 28891 28441 28903 28444
rect 28845 28435 28903 28441
rect 32401 28441 32413 28475
rect 32447 28472 32459 28475
rect 32447 28444 32628 28472
rect 32447 28441 32459 28444
rect 32401 28435 32459 28441
rect 23566 28404 23572 28416
rect 22388 28376 23572 28404
rect 21821 28367 21879 28373
rect 23566 28364 23572 28376
rect 23624 28364 23630 28416
rect 26326 28364 26332 28416
rect 26384 28404 26390 28416
rect 26605 28407 26663 28413
rect 26605 28404 26617 28407
rect 26384 28376 26617 28404
rect 26384 28364 26390 28376
rect 26605 28373 26617 28376
rect 26651 28373 26663 28407
rect 26605 28367 26663 28373
rect 27522 28364 27528 28416
rect 27580 28404 27586 28416
rect 27617 28407 27675 28413
rect 27617 28404 27629 28407
rect 27580 28376 27629 28404
rect 27580 28364 27586 28376
rect 27617 28373 27629 28376
rect 27663 28373 27675 28407
rect 27617 28367 27675 28373
rect 28994 28364 29000 28416
rect 29052 28404 29058 28416
rect 29641 28407 29699 28413
rect 29641 28404 29653 28407
rect 29052 28376 29653 28404
rect 29052 28364 29058 28376
rect 29641 28373 29653 28376
rect 29687 28373 29699 28407
rect 29641 28367 29699 28373
rect 30190 28364 30196 28416
rect 30248 28404 30254 28416
rect 32125 28407 32183 28413
rect 32125 28404 32137 28407
rect 30248 28376 32137 28404
rect 30248 28364 30254 28376
rect 32125 28373 32137 28376
rect 32171 28373 32183 28407
rect 32490 28404 32496 28416
rect 32451 28376 32496 28404
rect 32125 28367 32183 28373
rect 32490 28364 32496 28376
rect 32548 28364 32554 28416
rect 32600 28404 32628 28444
rect 32674 28432 32680 28484
rect 32732 28472 32738 28484
rect 33686 28481 33692 28484
rect 33663 28475 33692 28481
rect 32732 28444 32777 28472
rect 32732 28432 32738 28444
rect 33663 28441 33675 28475
rect 33663 28435 33692 28441
rect 33686 28432 33692 28435
rect 33744 28432 33750 28484
rect 33873 28475 33931 28481
rect 33873 28441 33885 28475
rect 33919 28472 33931 28475
rect 34054 28472 34060 28484
rect 33919 28444 34060 28472
rect 33919 28441 33931 28444
rect 33873 28435 33931 28441
rect 34054 28432 34060 28444
rect 34112 28472 34118 28484
rect 35544 28472 35572 28503
rect 34112 28444 35572 28472
rect 34112 28432 34118 28444
rect 32766 28404 32772 28416
rect 32600 28376 32772 28404
rect 32766 28364 32772 28376
rect 32824 28404 32830 28416
rect 34701 28407 34759 28413
rect 34701 28404 34713 28407
rect 32824 28376 34713 28404
rect 32824 28364 32830 28376
rect 34701 28373 34713 28376
rect 34747 28373 34759 28407
rect 34701 28367 34759 28373
rect 34790 28364 34796 28416
rect 34848 28404 34854 28416
rect 35636 28404 35664 28512
rect 35713 28509 35725 28512
rect 35759 28509 35771 28543
rect 35713 28503 35771 28509
rect 38102 28500 38108 28552
rect 38160 28540 38166 28552
rect 38160 28512 38205 28540
rect 38160 28500 38166 28512
rect 35710 28404 35716 28416
rect 34848 28376 35716 28404
rect 34848 28364 34854 28376
rect 35710 28364 35716 28376
rect 35768 28364 35774 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 8478 28200 8484 28212
rect 7300 28172 8484 28200
rect 7300 28076 7328 28172
rect 8478 28160 8484 28172
rect 8536 28200 8542 28212
rect 9858 28200 9864 28212
rect 8536 28172 9864 28200
rect 8536 28160 8542 28172
rect 9858 28160 9864 28172
rect 9916 28160 9922 28212
rect 10134 28160 10140 28212
rect 10192 28200 10198 28212
rect 10229 28203 10287 28209
rect 10229 28200 10241 28203
rect 10192 28172 10241 28200
rect 10192 28160 10198 28172
rect 10229 28169 10241 28172
rect 10275 28169 10287 28203
rect 10229 28163 10287 28169
rect 12406 28172 14228 28200
rect 7374 28092 7380 28144
rect 7432 28132 7438 28144
rect 12406 28132 12434 28172
rect 12802 28132 12808 28144
rect 7432 28104 8248 28132
rect 7432 28092 7438 28104
rect 6641 28067 6699 28073
rect 6641 28033 6653 28067
rect 6687 28064 6699 28067
rect 7282 28064 7288 28076
rect 6687 28036 7288 28064
rect 6687 28033 6699 28036
rect 6641 28027 6699 28033
rect 7282 28024 7288 28036
rect 7340 28024 7346 28076
rect 7742 28064 7748 28076
rect 7703 28036 7748 28064
rect 7742 28024 7748 28036
rect 7800 28024 7806 28076
rect 8021 28067 8079 28073
rect 8021 28033 8033 28067
rect 8067 28064 8079 28067
rect 8110 28064 8116 28076
rect 8067 28036 8116 28064
rect 8067 28033 8079 28036
rect 8021 28027 8079 28033
rect 8110 28024 8116 28036
rect 8168 28024 8174 28076
rect 8220 28073 8248 28104
rect 9416 28104 12434 28132
rect 12715 28104 12808 28132
rect 8205 28067 8263 28073
rect 8205 28033 8217 28067
rect 8251 28033 8263 28067
rect 8205 28027 8263 28033
rect 8220 27928 8248 28027
rect 8294 28024 8300 28076
rect 8352 28064 8358 28076
rect 9306 28064 9312 28076
rect 8352 28036 9312 28064
rect 8352 28024 8358 28036
rect 9306 28024 9312 28036
rect 9364 28024 9370 28076
rect 9416 28073 9444 28104
rect 12802 28092 12808 28104
rect 12860 28132 12866 28144
rect 13630 28132 13636 28144
rect 12860 28104 13636 28132
rect 12860 28092 12866 28104
rect 13630 28092 13636 28104
rect 13688 28092 13694 28144
rect 9401 28067 9459 28073
rect 9401 28033 9413 28067
rect 9447 28033 9459 28067
rect 9401 28027 9459 28033
rect 9858 28024 9864 28076
rect 9916 28064 9922 28076
rect 10137 28067 10195 28073
rect 10137 28064 10149 28067
rect 9916 28036 10149 28064
rect 9916 28024 9922 28036
rect 10137 28033 10149 28036
rect 10183 28064 10195 28067
rect 10226 28064 10232 28076
rect 10183 28036 10232 28064
rect 10183 28033 10195 28036
rect 10137 28027 10195 28033
rect 10226 28024 10232 28036
rect 10284 28024 10290 28076
rect 11698 28064 11704 28076
rect 11659 28036 11704 28064
rect 11698 28024 11704 28036
rect 11756 28024 11762 28076
rect 12529 28067 12587 28073
rect 12529 28064 12541 28067
rect 12406 28036 12541 28064
rect 9493 27999 9551 28005
rect 9493 27965 9505 27999
rect 9539 27965 9551 27999
rect 9493 27959 9551 27965
rect 9585 27999 9643 28005
rect 9585 27965 9597 27999
rect 9631 27996 9643 27999
rect 9674 27996 9680 28008
rect 9631 27968 9680 27996
rect 9631 27965 9643 27968
rect 9585 27959 9643 27965
rect 9508 27928 9536 27959
rect 9674 27956 9680 27968
rect 9732 27956 9738 28008
rect 11422 27956 11428 28008
rect 11480 27996 11486 28008
rect 11609 27999 11667 28005
rect 11609 27996 11621 27999
rect 11480 27968 11621 27996
rect 11480 27956 11486 27968
rect 11609 27965 11621 27968
rect 11655 27965 11667 27999
rect 11609 27959 11667 27965
rect 8220 27900 9536 27928
rect 6546 27860 6552 27872
rect 6507 27832 6552 27860
rect 6546 27820 6552 27832
rect 6604 27820 6610 27872
rect 7561 27863 7619 27869
rect 7561 27829 7573 27863
rect 7607 27860 7619 27863
rect 7834 27860 7840 27872
rect 7607 27832 7840 27860
rect 7607 27829 7619 27832
rect 7561 27823 7619 27829
rect 7834 27820 7840 27832
rect 7892 27820 7898 27872
rect 9122 27860 9128 27872
rect 9083 27832 9128 27860
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 9508 27860 9536 27900
rect 12069 27931 12127 27937
rect 12069 27897 12081 27931
rect 12115 27928 12127 27931
rect 12406 27928 12434 28036
rect 12529 28033 12541 28036
rect 12575 28033 12587 28067
rect 12710 28064 12716 28076
rect 12671 28036 12716 28064
rect 12529 28027 12587 28033
rect 12710 28024 12716 28036
rect 12768 28024 12774 28076
rect 12894 28024 12900 28076
rect 12952 28064 12958 28076
rect 13078 28064 13084 28076
rect 12952 28036 13084 28064
rect 12952 28024 12958 28036
rect 13078 28024 13084 28036
rect 13136 28024 13142 28076
rect 13538 28064 13544 28076
rect 13451 28036 13544 28064
rect 13538 28024 13544 28036
rect 13596 28024 13602 28076
rect 12618 27956 12624 28008
rect 12676 27996 12682 28008
rect 13556 27996 13584 28024
rect 12676 27968 13584 27996
rect 14200 27996 14228 28172
rect 14274 28160 14280 28212
rect 14332 28200 14338 28212
rect 14369 28203 14427 28209
rect 14369 28200 14381 28203
rect 14332 28172 14381 28200
rect 14332 28160 14338 28172
rect 14369 28169 14381 28172
rect 14415 28169 14427 28203
rect 14369 28163 14427 28169
rect 14458 28160 14464 28212
rect 14516 28200 14522 28212
rect 17310 28200 17316 28212
rect 14516 28172 17316 28200
rect 14516 28160 14522 28172
rect 15102 28141 15108 28144
rect 15089 28135 15108 28141
rect 15089 28101 15101 28135
rect 15089 28095 15108 28101
rect 15102 28092 15108 28095
rect 15160 28092 15166 28144
rect 15286 28132 15292 28144
rect 15247 28104 15292 28132
rect 15286 28092 15292 28104
rect 15344 28092 15350 28144
rect 15746 28092 15752 28144
rect 15804 28132 15810 28144
rect 15841 28135 15899 28141
rect 15841 28132 15853 28135
rect 15804 28104 15853 28132
rect 15804 28092 15810 28104
rect 15841 28101 15853 28104
rect 15887 28101 15899 28135
rect 15841 28095 15899 28101
rect 16684 28076 16712 28172
rect 17310 28160 17316 28172
rect 17368 28160 17374 28212
rect 17678 28160 17684 28212
rect 17736 28200 17742 28212
rect 18417 28203 18475 28209
rect 18417 28200 18429 28203
rect 17736 28172 18429 28200
rect 17736 28160 17742 28172
rect 18417 28169 18429 28172
rect 18463 28169 18475 28203
rect 18417 28163 18475 28169
rect 20349 28203 20407 28209
rect 20349 28169 20361 28203
rect 20395 28200 20407 28203
rect 20622 28200 20628 28212
rect 20395 28172 20628 28200
rect 20395 28169 20407 28172
rect 20349 28163 20407 28169
rect 20622 28160 20628 28172
rect 20680 28200 20686 28212
rect 21358 28200 21364 28212
rect 20680 28172 21364 28200
rect 20680 28160 20686 28172
rect 21358 28160 21364 28172
rect 21416 28160 21422 28212
rect 22002 28200 22008 28212
rect 21963 28172 22008 28200
rect 22002 28160 22008 28172
rect 22060 28160 22066 28212
rect 22646 28200 22652 28212
rect 22607 28172 22652 28200
rect 22646 28160 22652 28172
rect 22704 28160 22710 28212
rect 25866 28200 25872 28212
rect 25827 28172 25872 28200
rect 25866 28160 25872 28172
rect 25924 28160 25930 28212
rect 26973 28203 27031 28209
rect 26973 28169 26985 28203
rect 27019 28169 27031 28203
rect 29733 28203 29791 28209
rect 29733 28200 29745 28203
rect 26973 28163 27031 28169
rect 28092 28172 29745 28200
rect 16942 28132 16948 28144
rect 16903 28104 16948 28132
rect 16942 28092 16948 28104
rect 17000 28092 17006 28144
rect 18230 28132 18236 28144
rect 18170 28104 18236 28132
rect 18230 28092 18236 28104
rect 18288 28092 18294 28144
rect 21085 28135 21143 28141
rect 21085 28101 21097 28135
rect 21131 28132 21143 28135
rect 22922 28132 22928 28144
rect 21131 28104 22928 28132
rect 21131 28101 21143 28104
rect 21085 28095 21143 28101
rect 22922 28092 22928 28104
rect 22980 28092 22986 28144
rect 24857 28135 24915 28141
rect 24857 28101 24869 28135
rect 24903 28132 24915 28135
rect 26988 28132 27016 28163
rect 24903 28104 27016 28132
rect 27249 28135 27307 28141
rect 24903 28101 24915 28104
rect 24857 28095 24915 28101
rect 27249 28101 27261 28135
rect 27295 28132 27307 28135
rect 27430 28132 27436 28144
rect 27295 28104 27436 28132
rect 27295 28101 27307 28104
rect 27249 28095 27307 28101
rect 27430 28092 27436 28104
rect 27488 28132 27494 28144
rect 27890 28132 27896 28144
rect 27488 28104 27896 28132
rect 27488 28092 27494 28104
rect 27890 28092 27896 28104
rect 27948 28092 27954 28144
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28064 14519 28067
rect 14826 28064 14832 28076
rect 14507 28036 14832 28064
rect 14507 28033 14519 28036
rect 14461 28027 14519 28033
rect 14826 28024 14832 28036
rect 14884 28064 14890 28076
rect 15930 28064 15936 28076
rect 14884 28036 15936 28064
rect 14884 28024 14890 28036
rect 15930 28024 15936 28036
rect 15988 28024 15994 28076
rect 16666 28064 16672 28076
rect 16579 28036 16672 28064
rect 16666 28024 16672 28036
rect 16724 28024 16730 28076
rect 19061 28067 19119 28073
rect 19061 28033 19073 28067
rect 19107 28033 19119 28067
rect 19242 28064 19248 28076
rect 19203 28036 19248 28064
rect 19061 28027 19119 28033
rect 16942 27996 16948 28008
rect 14200 27968 16948 27996
rect 12676 27956 12682 27968
rect 12115 27900 12434 27928
rect 13556 27928 13584 27968
rect 16942 27956 16948 27968
rect 17000 27956 17006 28008
rect 17494 27956 17500 28008
rect 17552 27996 17558 28008
rect 19076 27996 19104 28027
rect 19242 28024 19248 28036
rect 19300 28024 19306 28076
rect 20165 28067 20223 28073
rect 20165 28033 20177 28067
rect 20211 28064 20223 28067
rect 20901 28067 20959 28073
rect 20901 28064 20913 28067
rect 20211 28036 20913 28064
rect 20211 28033 20223 28036
rect 20165 28027 20223 28033
rect 20901 28033 20913 28036
rect 20947 28033 20959 28067
rect 20901 28027 20959 28033
rect 22097 28067 22155 28073
rect 22097 28033 22109 28067
rect 22143 28064 22155 28067
rect 22186 28064 22192 28076
rect 22143 28036 22192 28064
rect 22143 28033 22155 28036
rect 22097 28027 22155 28033
rect 20180 27996 20208 28027
rect 22186 28024 22192 28036
rect 22244 28024 22250 28076
rect 22741 28067 22799 28073
rect 22741 28033 22753 28067
rect 22787 28064 22799 28067
rect 22830 28064 22836 28076
rect 22787 28036 22836 28064
rect 22787 28033 22799 28036
rect 22741 28027 22799 28033
rect 22830 28024 22836 28036
rect 22888 28024 22894 28076
rect 23750 28024 23756 28076
rect 23808 28024 23814 28076
rect 26050 28064 26056 28076
rect 26011 28036 26056 28064
rect 26050 28024 26056 28036
rect 26108 28024 26114 28076
rect 26326 28064 26332 28076
rect 26287 28036 26332 28064
rect 26326 28024 26332 28036
rect 26384 28024 26390 28076
rect 27154 28064 27160 28076
rect 27115 28036 27160 28064
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28033 27399 28067
rect 27522 28064 27528 28076
rect 27483 28036 27528 28064
rect 27341 28027 27399 28033
rect 17552 27968 19104 27996
rect 19168 27968 20208 27996
rect 22066 27968 25084 27996
rect 17552 27956 17558 27968
rect 19168 27928 19196 27968
rect 13556 27900 15332 27928
rect 12115 27897 12127 27900
rect 12069 27891 12127 27897
rect 9582 27860 9588 27872
rect 9508 27832 9588 27860
rect 9582 27820 9588 27832
rect 9640 27820 9646 27872
rect 12434 27820 12440 27872
rect 12492 27860 12498 27872
rect 12894 27860 12900 27872
rect 12492 27832 12900 27860
rect 12492 27820 12498 27832
rect 12894 27820 12900 27832
rect 12952 27820 12958 27872
rect 13078 27860 13084 27872
rect 13039 27832 13084 27860
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 13725 27863 13783 27869
rect 13725 27829 13737 27863
rect 13771 27860 13783 27863
rect 14826 27860 14832 27872
rect 13771 27832 14832 27860
rect 13771 27829 13783 27832
rect 13725 27823 13783 27829
rect 14826 27820 14832 27832
rect 14884 27820 14890 27872
rect 14918 27820 14924 27872
rect 14976 27860 14982 27872
rect 14976 27832 15021 27860
rect 14976 27820 14982 27832
rect 15102 27820 15108 27872
rect 15160 27860 15166 27872
rect 15304 27860 15332 27900
rect 17972 27900 19196 27928
rect 17972 27860 18000 27900
rect 19426 27888 19432 27940
rect 19484 27928 19490 27940
rect 22066 27928 22094 27968
rect 19484 27900 22094 27928
rect 19484 27888 19490 27900
rect 18874 27860 18880 27872
rect 15160 27832 15205 27860
rect 15304 27832 18000 27860
rect 18835 27832 18880 27860
rect 15160 27820 15166 27832
rect 18874 27820 18880 27832
rect 18932 27820 18938 27872
rect 21450 27820 21456 27872
rect 21508 27860 21514 27872
rect 21910 27860 21916 27872
rect 21508 27832 21916 27860
rect 21508 27820 21514 27832
rect 21910 27820 21916 27832
rect 21968 27820 21974 27872
rect 23385 27863 23443 27869
rect 23385 27829 23397 27863
rect 23431 27860 23443 27863
rect 23658 27860 23664 27872
rect 23431 27832 23664 27860
rect 23431 27829 23443 27832
rect 23385 27823 23443 27829
rect 23658 27820 23664 27832
rect 23716 27860 23722 27872
rect 24762 27860 24768 27872
rect 23716 27832 24768 27860
rect 23716 27820 23722 27832
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 25056 27860 25084 27968
rect 25130 27956 25136 28008
rect 25188 27996 25194 28008
rect 26234 27996 26240 28008
rect 25188 27968 25233 27996
rect 26195 27968 26240 27996
rect 25188 27956 25194 27968
rect 26234 27956 26240 27968
rect 26292 27996 26298 28008
rect 27356 27996 27384 28027
rect 27522 28024 27528 28036
rect 27580 28024 27586 28076
rect 26292 27968 27384 27996
rect 26292 27956 26298 27968
rect 25314 27888 25320 27940
rect 25372 27928 25378 27940
rect 26145 27931 26203 27937
rect 26145 27928 26157 27931
rect 25372 27900 26157 27928
rect 25372 27888 25378 27900
rect 26145 27897 26157 27900
rect 26191 27897 26203 27931
rect 26145 27891 26203 27897
rect 26878 27888 26884 27940
rect 26936 27928 26942 27940
rect 28092 27928 28120 28172
rect 29733 28169 29745 28172
rect 29779 28200 29791 28203
rect 30742 28200 30748 28212
rect 29779 28172 30748 28200
rect 29779 28169 29791 28172
rect 29733 28163 29791 28169
rect 30742 28160 30748 28172
rect 30800 28200 30806 28212
rect 30800 28172 31340 28200
rect 30800 28160 30806 28172
rect 29822 28132 29828 28144
rect 28920 28104 29828 28132
rect 28920 28073 28948 28104
rect 29822 28092 29828 28104
rect 29880 28092 29886 28144
rect 28169 28067 28227 28073
rect 28169 28033 28181 28067
rect 28215 28064 28227 28067
rect 28905 28067 28963 28073
rect 28905 28064 28917 28067
rect 28215 28036 28917 28064
rect 28215 28033 28227 28036
rect 28169 28027 28227 28033
rect 28905 28033 28917 28036
rect 28951 28033 28963 28067
rect 28905 28027 28963 28033
rect 26936 27900 28120 27928
rect 26936 27888 26942 27900
rect 28184 27860 28212 28027
rect 28994 28024 29000 28076
rect 29052 28064 29058 28076
rect 29641 28067 29699 28073
rect 29641 28064 29653 28067
rect 29052 28036 29653 28064
rect 29052 28024 29058 28036
rect 29641 28033 29653 28036
rect 29687 28033 29699 28067
rect 30374 28064 30380 28076
rect 30287 28036 30380 28064
rect 29641 28027 29699 28033
rect 30374 28024 30380 28036
rect 30432 28024 30438 28076
rect 31312 28073 31340 28172
rect 32122 28160 32128 28212
rect 32180 28200 32186 28212
rect 32766 28209 32772 28212
rect 32585 28203 32643 28209
rect 32585 28200 32597 28203
rect 32180 28172 32597 28200
rect 32180 28160 32186 28172
rect 32585 28169 32597 28172
rect 32631 28169 32643 28203
rect 32585 28163 32643 28169
rect 32753 28203 32772 28209
rect 32753 28169 32765 28203
rect 32753 28163 32772 28169
rect 32766 28160 32772 28163
rect 32824 28160 32830 28212
rect 34882 28200 34888 28212
rect 33796 28172 34888 28200
rect 32950 28132 32956 28144
rect 32911 28104 32956 28132
rect 32950 28092 32956 28104
rect 33008 28092 33014 28144
rect 33686 28132 33692 28144
rect 33060 28104 33692 28132
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28064 31355 28067
rect 31386 28064 31392 28076
rect 31343 28036 31392 28064
rect 31343 28033 31355 28036
rect 31297 28027 31355 28033
rect 31386 28024 31392 28036
rect 31444 28024 31450 28076
rect 31478 28024 31484 28076
rect 31536 28064 31542 28076
rect 33060 28064 33088 28104
rect 33686 28092 33692 28104
rect 33744 28092 33750 28144
rect 33796 28141 33824 28172
rect 34882 28160 34888 28172
rect 34940 28160 34946 28212
rect 34974 28160 34980 28212
rect 35032 28200 35038 28212
rect 36265 28203 36323 28209
rect 36265 28200 36277 28203
rect 35032 28172 36277 28200
rect 35032 28160 35038 28172
rect 36265 28169 36277 28172
rect 36311 28169 36323 28203
rect 36265 28163 36323 28169
rect 33781 28135 33839 28141
rect 33781 28101 33793 28135
rect 33827 28101 33839 28135
rect 33781 28095 33839 28101
rect 34057 28135 34115 28141
rect 34057 28101 34069 28135
rect 34103 28132 34115 28135
rect 34793 28135 34851 28141
rect 34793 28132 34805 28135
rect 34103 28104 34805 28132
rect 34103 28101 34115 28104
rect 34057 28095 34115 28101
rect 34793 28101 34805 28104
rect 34839 28101 34851 28135
rect 34793 28095 34851 28101
rect 31536 28036 33088 28064
rect 31536 28024 31542 28036
rect 33134 28024 33140 28076
rect 33192 28064 33198 28076
rect 33594 28073 33600 28076
rect 33551 28067 33600 28073
rect 33551 28064 33563 28067
rect 33192 28036 33563 28064
rect 33192 28024 33198 28036
rect 33551 28033 33563 28036
rect 33597 28033 33600 28067
rect 33551 28027 33600 28033
rect 33594 28024 33600 28027
rect 33652 28064 33658 28076
rect 33873 28067 33931 28073
rect 33652 28036 33699 28064
rect 33652 28024 33658 28036
rect 33873 28033 33885 28067
rect 33919 28033 33931 28067
rect 33873 28027 33931 28033
rect 29086 27996 29092 28008
rect 28999 27968 29092 27996
rect 29086 27956 29092 27968
rect 29144 27996 29150 28008
rect 30006 27996 30012 28008
rect 29144 27968 30012 27996
rect 29144 27956 29150 27968
rect 30006 27956 30012 27968
rect 30064 27956 30070 28008
rect 30392 27996 30420 28024
rect 31662 27996 31668 28008
rect 30392 27968 31668 27996
rect 31662 27956 31668 27968
rect 31720 27956 31726 28008
rect 33318 27956 33324 28008
rect 33376 27996 33382 28008
rect 33413 27999 33471 28005
rect 33413 27996 33425 27999
rect 33376 27968 33425 27996
rect 33376 27956 33382 27968
rect 33413 27965 33425 27968
rect 33459 27965 33471 27999
rect 33413 27959 33471 27965
rect 28353 27931 28411 27937
rect 28353 27897 28365 27931
rect 28399 27928 28411 27931
rect 28718 27928 28724 27940
rect 28399 27900 28724 27928
rect 28399 27897 28411 27900
rect 28353 27891 28411 27897
rect 28718 27888 28724 27900
rect 28776 27928 28782 27940
rect 30650 27928 30656 27940
rect 28776 27900 30656 27928
rect 28776 27888 28782 27900
rect 30650 27888 30656 27900
rect 30708 27888 30714 27940
rect 31570 27928 31576 27940
rect 30944 27900 31576 27928
rect 30944 27872 30972 27900
rect 31570 27888 31576 27900
rect 31628 27888 31634 27940
rect 32490 27888 32496 27940
rect 32548 27928 32554 27940
rect 32548 27900 32812 27928
rect 32548 27888 32554 27900
rect 25056 27832 28212 27860
rect 30469 27863 30527 27869
rect 30469 27829 30481 27863
rect 30515 27860 30527 27863
rect 30926 27860 30932 27872
rect 30515 27832 30932 27860
rect 30515 27829 30527 27832
rect 30469 27823 30527 27829
rect 30926 27820 30932 27832
rect 30984 27820 30990 27872
rect 31478 27860 31484 27872
rect 31439 27832 31484 27860
rect 31478 27820 31484 27832
rect 31536 27820 31542 27872
rect 32784 27869 32812 27900
rect 32769 27863 32827 27869
rect 32769 27829 32781 27863
rect 32815 27860 32827 27863
rect 33502 27860 33508 27872
rect 32815 27832 33508 27860
rect 32815 27829 32827 27832
rect 32769 27823 32827 27829
rect 33502 27820 33508 27832
rect 33560 27820 33566 27872
rect 33888 27860 33916 28027
rect 35894 28024 35900 28076
rect 35952 28024 35958 28076
rect 37829 28067 37887 28073
rect 37829 28033 37841 28067
rect 37875 28064 37887 28067
rect 38102 28064 38108 28076
rect 37875 28036 38108 28064
rect 37875 28033 37887 28036
rect 37829 28027 37887 28033
rect 38102 28024 38108 28036
rect 38160 28024 38166 28076
rect 34514 27996 34520 28008
rect 34475 27968 34520 27996
rect 34514 27956 34520 27968
rect 34572 27956 34578 28008
rect 34606 27860 34612 27872
rect 33888 27832 34612 27860
rect 34606 27820 34612 27832
rect 34664 27820 34670 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 6567 27659 6625 27665
rect 6567 27625 6579 27659
rect 6613 27656 6625 27659
rect 7285 27659 7343 27665
rect 7285 27656 7297 27659
rect 6613 27628 7297 27656
rect 6613 27625 6625 27628
rect 6567 27619 6625 27625
rect 7285 27625 7297 27628
rect 7331 27625 7343 27659
rect 7285 27619 7343 27625
rect 11698 27616 11704 27668
rect 11756 27656 11762 27668
rect 11793 27659 11851 27665
rect 11793 27656 11805 27659
rect 11756 27628 11805 27656
rect 11756 27616 11762 27628
rect 11793 27625 11805 27628
rect 11839 27656 11851 27659
rect 12802 27656 12808 27668
rect 11839 27628 12808 27656
rect 11839 27625 11851 27628
rect 11793 27619 11851 27625
rect 12802 27616 12808 27628
rect 12860 27616 12866 27668
rect 13078 27616 13084 27668
rect 13136 27656 13142 27668
rect 13277 27659 13335 27665
rect 13277 27656 13289 27659
rect 13136 27628 13289 27656
rect 13136 27616 13142 27628
rect 13277 27625 13289 27628
rect 13323 27625 13335 27659
rect 16669 27659 16727 27665
rect 13277 27619 13335 27625
rect 14844 27628 15056 27656
rect 7006 27548 7012 27600
rect 7064 27588 7070 27600
rect 12250 27588 12256 27600
rect 7064 27560 12256 27588
rect 7064 27548 7070 27560
rect 6178 27480 6184 27532
rect 6236 27520 6242 27532
rect 6825 27523 6883 27529
rect 6825 27520 6837 27523
rect 6236 27492 6837 27520
rect 6236 27480 6242 27492
rect 6825 27489 6837 27492
rect 6871 27489 6883 27523
rect 6825 27483 6883 27489
rect 7484 27461 7512 27560
rect 12250 27548 12256 27560
rect 12308 27548 12314 27600
rect 14458 27548 14464 27600
rect 14516 27588 14522 27600
rect 14844 27588 14872 27628
rect 14516 27560 14872 27588
rect 14516 27548 14522 27560
rect 14918 27548 14924 27600
rect 14976 27548 14982 27600
rect 15028 27588 15056 27628
rect 16669 27625 16681 27659
rect 16715 27656 16727 27659
rect 16758 27656 16764 27668
rect 16715 27628 16764 27656
rect 16715 27625 16727 27628
rect 16669 27619 16727 27625
rect 16758 27616 16764 27628
rect 16816 27616 16822 27668
rect 17402 27616 17408 27668
rect 17460 27656 17466 27668
rect 17589 27659 17647 27665
rect 17589 27656 17601 27659
rect 17460 27628 17601 27656
rect 17460 27616 17466 27628
rect 17589 27625 17601 27628
rect 17635 27625 17647 27659
rect 19242 27656 19248 27668
rect 17589 27619 17647 27625
rect 17972 27628 18276 27656
rect 19203 27628 19248 27656
rect 16850 27588 16856 27600
rect 15028 27560 16856 27588
rect 16850 27548 16856 27560
rect 16908 27588 16914 27600
rect 17972 27588 18000 27628
rect 16908 27560 18000 27588
rect 18049 27591 18107 27597
rect 16908 27548 16914 27560
rect 18049 27557 18061 27591
rect 18095 27588 18107 27591
rect 18138 27588 18144 27600
rect 18095 27560 18144 27588
rect 18095 27557 18107 27560
rect 18049 27551 18107 27557
rect 18138 27548 18144 27560
rect 18196 27548 18202 27600
rect 18248 27588 18276 27628
rect 19242 27616 19248 27628
rect 19300 27616 19306 27668
rect 21910 27616 21916 27668
rect 21968 27656 21974 27668
rect 28166 27656 28172 27668
rect 21968 27628 28172 27656
rect 21968 27616 21974 27628
rect 28166 27616 28172 27628
rect 28224 27616 28230 27668
rect 28353 27659 28411 27665
rect 28353 27625 28365 27659
rect 28399 27625 28411 27659
rect 28353 27619 28411 27625
rect 22278 27588 22284 27600
rect 18248 27560 22284 27588
rect 22278 27548 22284 27560
rect 22336 27548 22342 27600
rect 23750 27588 23756 27600
rect 23711 27560 23756 27588
rect 23750 27548 23756 27560
rect 23808 27548 23814 27600
rect 24489 27591 24547 27597
rect 24489 27557 24501 27591
rect 24535 27588 24547 27591
rect 27338 27588 27344 27600
rect 24535 27560 27344 27588
rect 24535 27557 24547 27560
rect 24489 27551 24547 27557
rect 9582 27520 9588 27532
rect 9543 27492 9588 27520
rect 9582 27480 9588 27492
rect 9640 27480 9646 27532
rect 9674 27480 9680 27532
rect 9732 27520 9738 27532
rect 9732 27492 9777 27520
rect 9732 27480 9738 27492
rect 9950 27480 9956 27532
rect 10008 27520 10014 27532
rect 10965 27523 11023 27529
rect 10965 27520 10977 27523
rect 10008 27492 10977 27520
rect 10008 27480 10014 27492
rect 10965 27489 10977 27492
rect 11011 27489 11023 27523
rect 12710 27520 12716 27532
rect 10965 27483 11023 27489
rect 11992 27492 12716 27520
rect 7469 27455 7527 27461
rect 7469 27421 7481 27455
rect 7515 27421 7527 27455
rect 7834 27452 7840 27464
rect 7795 27424 7840 27452
rect 7469 27415 7527 27421
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 9306 27412 9312 27464
rect 9364 27452 9370 27464
rect 9493 27455 9551 27461
rect 9493 27452 9505 27455
rect 9364 27424 9505 27452
rect 9364 27412 9370 27424
rect 9493 27421 9505 27424
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 9769 27455 9827 27461
rect 9769 27421 9781 27455
rect 9815 27452 9827 27455
rect 10870 27452 10876 27464
rect 9815 27424 10876 27452
rect 9815 27421 9827 27424
rect 9769 27415 9827 27421
rect 10870 27412 10876 27424
rect 10928 27412 10934 27464
rect 11057 27455 11115 27461
rect 11057 27421 11069 27455
rect 11103 27452 11115 27455
rect 11882 27452 11888 27464
rect 11103 27424 11888 27452
rect 11103 27421 11115 27424
rect 11057 27415 11115 27421
rect 11882 27412 11888 27424
rect 11940 27412 11946 27464
rect 6546 27384 6552 27396
rect 6118 27356 6552 27384
rect 6546 27344 6552 27356
rect 6604 27344 6610 27396
rect 7374 27344 7380 27396
rect 7432 27384 7438 27396
rect 7561 27387 7619 27393
rect 7561 27384 7573 27387
rect 7432 27356 7573 27384
rect 7432 27344 7438 27356
rect 7561 27353 7573 27356
rect 7607 27353 7619 27387
rect 7561 27347 7619 27353
rect 7653 27387 7711 27393
rect 7653 27353 7665 27387
rect 7699 27384 7711 27387
rect 8018 27384 8024 27396
rect 7699 27356 8024 27384
rect 7699 27353 7711 27356
rect 7653 27347 7711 27353
rect 8018 27344 8024 27356
rect 8076 27384 8082 27396
rect 11992 27384 12020 27492
rect 12710 27480 12716 27492
rect 12768 27480 12774 27532
rect 14826 27480 14832 27532
rect 14884 27480 14890 27532
rect 14936 27520 14964 27548
rect 14936 27492 15608 27520
rect 13538 27412 13544 27464
rect 13596 27452 13602 27464
rect 14277 27455 14335 27461
rect 13596 27424 13641 27452
rect 13596 27412 13602 27424
rect 14277 27421 14289 27455
rect 14323 27452 14335 27455
rect 14734 27452 14740 27464
rect 14323 27424 14740 27452
rect 14323 27421 14335 27424
rect 14277 27415 14335 27421
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 14844 27452 14872 27480
rect 15580 27461 15608 27492
rect 16114 27480 16120 27532
rect 16172 27520 16178 27532
rect 17681 27523 17739 27529
rect 17681 27520 17693 27523
rect 16172 27492 17693 27520
rect 16172 27480 16178 27492
rect 17681 27489 17693 27492
rect 17727 27520 17739 27523
rect 18598 27520 18604 27532
rect 17727 27492 18604 27520
rect 17727 27489 17739 27492
rect 17681 27483 17739 27489
rect 18598 27480 18604 27492
rect 18656 27480 18662 27532
rect 19613 27523 19671 27529
rect 19613 27489 19625 27523
rect 19659 27520 19671 27523
rect 20257 27523 20315 27529
rect 20257 27520 20269 27523
rect 19659 27492 20269 27520
rect 19659 27489 19671 27492
rect 19613 27483 19671 27489
rect 20257 27489 20269 27492
rect 20303 27489 20315 27523
rect 20257 27483 20315 27489
rect 14921 27455 14979 27461
rect 14921 27452 14933 27455
rect 14844 27424 14933 27452
rect 14921 27421 14933 27424
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27421 15531 27455
rect 15473 27415 15531 27421
rect 15565 27455 15623 27461
rect 15565 27421 15577 27455
rect 15611 27421 15623 27455
rect 16206 27452 16212 27464
rect 16167 27424 16212 27452
rect 15565 27415 15623 27421
rect 14829 27387 14887 27393
rect 14829 27384 14841 27387
rect 8076 27356 12020 27384
rect 12834 27356 14841 27384
rect 8076 27344 8082 27356
rect 14829 27353 14841 27356
rect 14875 27353 14887 27387
rect 15488 27384 15516 27415
rect 16206 27412 16212 27424
rect 16264 27412 16270 27464
rect 16301 27455 16359 27461
rect 16301 27421 16313 27455
rect 16347 27452 16359 27455
rect 16390 27452 16396 27464
rect 16347 27424 16396 27452
rect 16347 27421 16359 27424
rect 16301 27415 16359 27421
rect 16390 27412 16396 27424
rect 16448 27412 16454 27464
rect 16485 27455 16543 27461
rect 16485 27421 16497 27455
rect 16531 27452 16543 27455
rect 17402 27452 17408 27464
rect 16531 27424 17408 27452
rect 16531 27421 16543 27424
rect 16485 27415 16543 27421
rect 17402 27412 17408 27424
rect 17460 27412 17466 27464
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 18322 27452 18328 27464
rect 17911 27424 18328 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 18322 27412 18328 27424
rect 18380 27412 18386 27464
rect 18414 27412 18420 27464
rect 18472 27452 18478 27464
rect 18509 27455 18567 27461
rect 18509 27452 18521 27455
rect 18472 27424 18521 27452
rect 18472 27412 18478 27424
rect 18509 27421 18521 27424
rect 18555 27448 18567 27455
rect 19426 27452 19432 27464
rect 18555 27421 18644 27448
rect 19387 27424 19432 27452
rect 18509 27420 18644 27421
rect 18509 27415 18567 27420
rect 15654 27384 15660 27396
rect 15488 27356 15660 27384
rect 14829 27347 14887 27353
rect 15654 27344 15660 27356
rect 15712 27384 15718 27396
rect 17589 27387 17647 27393
rect 17589 27384 17601 27387
rect 15712 27356 17601 27384
rect 15712 27344 15718 27356
rect 17589 27353 17601 27356
rect 17635 27353 17647 27387
rect 18616 27384 18644 27420
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 20349 27455 20407 27461
rect 20349 27421 20361 27455
rect 20395 27452 20407 27455
rect 20438 27452 20444 27464
rect 20395 27424 20444 27452
rect 20395 27421 20407 27424
rect 20349 27415 20407 27421
rect 19720 27384 19748 27415
rect 18616 27356 19748 27384
rect 17589 27347 17647 27353
rect 5077 27319 5135 27325
rect 5077 27285 5089 27319
rect 5123 27316 5135 27319
rect 7098 27316 7104 27328
rect 5123 27288 7104 27316
rect 5123 27285 5135 27288
rect 5077 27279 5135 27285
rect 7098 27276 7104 27288
rect 7156 27276 7162 27328
rect 9306 27316 9312 27328
rect 9267 27288 9312 27316
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 14090 27316 14096 27328
rect 14051 27288 14096 27316
rect 14090 27276 14096 27288
rect 14148 27276 14154 27328
rect 15749 27319 15807 27325
rect 15749 27285 15761 27319
rect 15795 27316 15807 27319
rect 16206 27316 16212 27328
rect 15795 27288 16212 27316
rect 15795 27285 15807 27288
rect 15749 27279 15807 27285
rect 16206 27276 16212 27288
rect 16264 27276 16270 27328
rect 18601 27319 18659 27325
rect 18601 27285 18613 27319
rect 18647 27316 18659 27319
rect 18690 27316 18696 27328
rect 18647 27288 18696 27316
rect 18647 27285 18659 27288
rect 18601 27279 18659 27285
rect 18690 27276 18696 27288
rect 18748 27276 18754 27328
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 20180 27316 20208 27415
rect 20438 27412 20444 27424
rect 20496 27412 20502 27464
rect 20622 27412 20628 27464
rect 20680 27452 20686 27464
rect 20993 27455 21051 27461
rect 20993 27452 21005 27455
rect 20680 27424 21005 27452
rect 20680 27412 20686 27424
rect 20993 27421 21005 27424
rect 21039 27421 21051 27455
rect 20993 27415 21051 27421
rect 22649 27455 22707 27461
rect 22649 27421 22661 27455
rect 22695 27452 22707 27455
rect 23474 27452 23480 27464
rect 22695 27424 23480 27452
rect 22695 27421 22707 27424
rect 22649 27415 22707 27421
rect 23474 27412 23480 27424
rect 23532 27412 23538 27464
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 23661 27455 23719 27461
rect 23661 27452 23673 27455
rect 23624 27424 23673 27452
rect 23624 27412 23630 27424
rect 23661 27421 23673 27424
rect 23707 27452 23719 27455
rect 24504 27452 24532 27551
rect 27338 27548 27344 27560
rect 27396 27548 27402 27600
rect 27522 27548 27528 27600
rect 27580 27588 27586 27600
rect 28368 27588 28396 27619
rect 28442 27616 28448 27668
rect 28500 27656 28506 27668
rect 31110 27656 31116 27668
rect 28500 27628 31116 27656
rect 28500 27616 28506 27628
rect 31110 27616 31116 27628
rect 31168 27656 31174 27668
rect 31478 27656 31484 27668
rect 31168 27628 31484 27656
rect 31168 27616 31174 27628
rect 31478 27616 31484 27628
rect 31536 27616 31542 27668
rect 32950 27616 32956 27668
rect 33008 27656 33014 27668
rect 33965 27659 34023 27665
rect 33965 27656 33977 27659
rect 33008 27628 33977 27656
rect 33008 27616 33014 27628
rect 33965 27625 33977 27628
rect 34011 27656 34023 27659
rect 34011 27628 34836 27656
rect 34011 27625 34023 27628
rect 33965 27619 34023 27625
rect 27580 27560 28396 27588
rect 28629 27591 28687 27597
rect 27580 27548 27586 27560
rect 28629 27557 28641 27591
rect 28675 27588 28687 27591
rect 28810 27588 28816 27600
rect 28675 27560 28816 27588
rect 28675 27557 28687 27560
rect 28629 27551 28687 27557
rect 28810 27548 28816 27560
rect 28868 27548 28874 27600
rect 30742 27588 30748 27600
rect 30300 27560 30748 27588
rect 25593 27523 25651 27529
rect 25593 27489 25605 27523
rect 25639 27520 25651 27523
rect 26421 27523 26479 27529
rect 26421 27520 26433 27523
rect 25639 27492 26433 27520
rect 25639 27489 25651 27492
rect 25593 27483 25651 27489
rect 26421 27489 26433 27492
rect 26467 27489 26479 27523
rect 26421 27483 26479 27489
rect 26513 27523 26571 27529
rect 26513 27489 26525 27523
rect 26559 27520 26571 27523
rect 28074 27520 28080 27532
rect 26559 27492 28080 27520
rect 26559 27489 26571 27492
rect 26513 27483 26571 27489
rect 24670 27452 24676 27464
rect 23707 27424 24532 27452
rect 24631 27424 24676 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 24670 27412 24676 27424
rect 24728 27412 24734 27464
rect 25682 27452 25688 27464
rect 25643 27424 25688 27452
rect 25682 27412 25688 27424
rect 25740 27412 25746 27464
rect 26050 27412 26056 27464
rect 26108 27452 26114 27464
rect 26326 27452 26332 27464
rect 26108 27424 26332 27452
rect 26108 27412 26114 27424
rect 26326 27412 26332 27424
rect 26384 27412 26390 27464
rect 26605 27455 26663 27461
rect 26605 27421 26617 27455
rect 26651 27452 26663 27455
rect 26786 27452 26792 27464
rect 26651 27424 26792 27452
rect 26651 27421 26663 27424
rect 26605 27415 26663 27421
rect 26786 27412 26792 27424
rect 26844 27412 26850 27464
rect 26970 27412 26976 27464
rect 27028 27452 27034 27464
rect 27356 27461 27384 27492
rect 28074 27480 28080 27492
rect 28132 27480 28138 27532
rect 28166 27480 28172 27532
rect 28224 27520 28230 27532
rect 28224 27492 29592 27520
rect 28224 27480 28230 27492
rect 27157 27455 27215 27461
rect 27157 27452 27169 27455
rect 27028 27424 27169 27452
rect 27028 27412 27034 27424
rect 27157 27421 27169 27424
rect 27203 27421 27215 27455
rect 27157 27415 27215 27421
rect 27341 27455 27399 27461
rect 27341 27421 27353 27455
rect 27387 27421 27399 27455
rect 27522 27452 27528 27464
rect 27483 27424 27528 27452
rect 27341 27415 27399 27421
rect 27522 27412 27528 27424
rect 27580 27412 27586 27464
rect 27706 27412 27712 27464
rect 27764 27412 27770 27464
rect 27798 27412 27804 27464
rect 27856 27452 27862 27464
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 27856 27424 28365 27452
rect 27856 27412 27862 27424
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 28353 27415 28411 27421
rect 28442 27412 28448 27464
rect 28500 27452 28506 27464
rect 29564 27461 29592 27492
rect 29549 27455 29607 27461
rect 28500 27424 28545 27452
rect 28500 27412 28506 27424
rect 29549 27421 29561 27455
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 30193 27455 30251 27461
rect 30193 27421 30205 27455
rect 30239 27452 30251 27455
rect 30300 27452 30328 27560
rect 30742 27548 30748 27560
rect 30800 27588 30806 27600
rect 30800 27560 31524 27588
rect 30800 27548 30806 27560
rect 31110 27520 31116 27532
rect 30484 27492 31116 27520
rect 30484 27461 30512 27492
rect 31110 27480 31116 27492
rect 31168 27520 31174 27532
rect 31496 27529 31524 27560
rect 34606 27548 34612 27600
rect 34664 27588 34670 27600
rect 34701 27591 34759 27597
rect 34701 27588 34713 27591
rect 34664 27560 34713 27588
rect 34664 27548 34670 27560
rect 34701 27557 34713 27560
rect 34747 27557 34759 27591
rect 34808 27588 34836 27628
rect 34808 27560 35296 27588
rect 34701 27551 34759 27557
rect 31297 27523 31355 27529
rect 31297 27520 31309 27523
rect 31168 27492 31309 27520
rect 31168 27480 31174 27492
rect 31297 27489 31309 27492
rect 31343 27489 31355 27523
rect 31297 27483 31355 27489
rect 31481 27523 31539 27529
rect 31481 27489 31493 27523
rect 31527 27489 31539 27523
rect 31481 27483 31539 27489
rect 32309 27523 32367 27529
rect 32309 27489 32321 27523
rect 32355 27520 32367 27523
rect 32674 27520 32680 27532
rect 32355 27492 32680 27520
rect 32355 27489 32367 27492
rect 32309 27483 32367 27489
rect 32674 27480 32680 27492
rect 32732 27480 32738 27532
rect 33502 27480 33508 27532
rect 33560 27520 33566 27532
rect 34422 27520 34428 27532
rect 33560 27492 34428 27520
rect 33560 27480 33566 27492
rect 34422 27480 34428 27492
rect 34480 27520 34486 27532
rect 34480 27492 35204 27520
rect 34480 27480 34486 27492
rect 30239 27424 30328 27452
rect 30469 27455 30527 27461
rect 30239 27421 30251 27424
rect 30193 27415 30251 27421
rect 30469 27421 30481 27455
rect 30515 27421 30527 27455
rect 31202 27452 31208 27464
rect 31163 27424 31208 27452
rect 30469 27415 30527 27421
rect 31202 27412 31208 27424
rect 31260 27412 31266 27464
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27421 31447 27455
rect 32582 27452 32588 27464
rect 32543 27424 32588 27452
rect 31389 27415 31447 27421
rect 23492 27384 23520 27412
rect 24578 27384 24584 27396
rect 23492 27356 24584 27384
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 27430 27384 27436 27396
rect 27391 27356 27436 27384
rect 27430 27344 27436 27356
rect 27488 27344 27494 27396
rect 19116 27288 20208 27316
rect 19116 27276 19122 27288
rect 20346 27276 20352 27328
rect 20404 27316 20410 27328
rect 20901 27319 20959 27325
rect 20901 27316 20913 27319
rect 20404 27288 20913 27316
rect 20404 27276 20410 27288
rect 20901 27285 20913 27288
rect 20947 27285 20959 27319
rect 22738 27316 22744 27328
rect 22699 27288 22744 27316
rect 20901 27279 20959 27285
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 24670 27276 24676 27328
rect 24728 27316 24734 27328
rect 27724 27325 27752 27412
rect 28169 27387 28227 27393
rect 28169 27353 28181 27387
rect 28215 27384 28227 27387
rect 29730 27384 29736 27396
rect 28215 27356 29736 27384
rect 28215 27353 28227 27356
rect 28169 27347 28227 27353
rect 29730 27344 29736 27356
rect 29788 27344 29794 27396
rect 30285 27387 30343 27393
rect 30285 27353 30297 27387
rect 30331 27384 30343 27387
rect 30374 27384 30380 27396
rect 30331 27356 30380 27384
rect 30331 27353 30343 27356
rect 30285 27347 30343 27353
rect 30374 27344 30380 27356
rect 30432 27384 30438 27396
rect 31404 27384 31432 27415
rect 32582 27412 32588 27424
rect 32640 27452 32646 27464
rect 32950 27452 32956 27464
rect 32640 27424 32956 27452
rect 32640 27412 32646 27424
rect 32950 27412 32956 27424
rect 33008 27412 33014 27464
rect 35176 27461 35204 27492
rect 34885 27455 34943 27461
rect 34885 27421 34897 27455
rect 34931 27421 34943 27455
rect 34885 27415 34943 27421
rect 35161 27455 35219 27461
rect 35161 27421 35173 27455
rect 35207 27421 35219 27455
rect 35161 27415 35219 27421
rect 30432 27356 31432 27384
rect 30432 27344 30438 27356
rect 33594 27344 33600 27396
rect 33652 27384 33658 27396
rect 33781 27387 33839 27393
rect 33781 27384 33793 27387
rect 33652 27356 33793 27384
rect 33652 27344 33658 27356
rect 33781 27353 33793 27356
rect 33827 27384 33839 27387
rect 34900 27384 34928 27415
rect 33827 27356 34928 27384
rect 35069 27387 35127 27393
rect 33827 27353 33839 27356
rect 33781 27347 33839 27353
rect 35069 27353 35081 27387
rect 35115 27384 35127 27387
rect 35268 27384 35296 27560
rect 38105 27523 38163 27529
rect 38105 27489 38117 27523
rect 38151 27520 38163 27523
rect 38654 27520 38660 27532
rect 38151 27492 38660 27520
rect 38151 27489 38163 27492
rect 38105 27483 38163 27489
rect 38654 27480 38660 27492
rect 38712 27480 38718 27532
rect 36262 27452 36268 27464
rect 36223 27424 36268 27452
rect 36262 27412 36268 27424
rect 36320 27412 36326 27464
rect 35526 27384 35532 27396
rect 35115 27356 35532 27384
rect 35115 27353 35127 27356
rect 35069 27347 35127 27353
rect 35526 27344 35532 27356
rect 35584 27344 35590 27396
rect 36449 27387 36507 27393
rect 36449 27353 36461 27387
rect 36495 27384 36507 27387
rect 37366 27384 37372 27396
rect 36495 27356 37372 27384
rect 36495 27353 36507 27356
rect 36449 27347 36507 27353
rect 37366 27344 37372 27356
rect 37424 27344 37430 27396
rect 26145 27319 26203 27325
rect 26145 27316 26157 27319
rect 24728 27288 26157 27316
rect 24728 27276 24734 27288
rect 26145 27285 26157 27288
rect 26191 27285 26203 27319
rect 26145 27279 26203 27285
rect 27709 27319 27767 27325
rect 27709 27285 27721 27319
rect 27755 27285 27767 27319
rect 27709 27279 27767 27285
rect 27890 27276 27896 27328
rect 27948 27316 27954 27328
rect 29086 27316 29092 27328
rect 27948 27288 29092 27316
rect 27948 27276 27954 27288
rect 29086 27276 29092 27288
rect 29144 27276 29150 27328
rect 29546 27276 29552 27328
rect 29604 27316 29610 27328
rect 29641 27319 29699 27325
rect 29641 27316 29653 27319
rect 29604 27288 29653 27316
rect 29604 27276 29610 27288
rect 29641 27285 29653 27288
rect 29687 27285 29699 27319
rect 29641 27279 29699 27285
rect 30558 27276 30564 27328
rect 30616 27316 30622 27328
rect 30653 27319 30711 27325
rect 30653 27316 30665 27319
rect 30616 27288 30665 27316
rect 30616 27276 30622 27288
rect 30653 27285 30665 27288
rect 30699 27285 30711 27319
rect 30653 27279 30711 27285
rect 31665 27319 31723 27325
rect 31665 27285 31677 27319
rect 31711 27316 31723 27319
rect 32122 27316 32128 27328
rect 31711 27288 32128 27316
rect 31711 27285 31723 27288
rect 31665 27279 31723 27285
rect 32122 27276 32128 27288
rect 32180 27276 32186 27328
rect 33502 27276 33508 27328
rect 33560 27316 33566 27328
rect 33981 27319 34039 27325
rect 33981 27316 33993 27319
rect 33560 27288 33993 27316
rect 33560 27276 33566 27288
rect 33981 27285 33993 27288
rect 34027 27285 34039 27319
rect 33981 27279 34039 27285
rect 34149 27319 34207 27325
rect 34149 27285 34161 27319
rect 34195 27316 34207 27319
rect 34698 27316 34704 27328
rect 34195 27288 34704 27316
rect 34195 27285 34207 27288
rect 34149 27279 34207 27285
rect 34698 27276 34704 27288
rect 34756 27276 34762 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 8849 27115 8907 27121
rect 8849 27081 8861 27115
rect 8895 27112 8907 27115
rect 9674 27112 9680 27124
rect 8895 27084 9680 27112
rect 8895 27081 8907 27084
rect 8849 27075 8907 27081
rect 9674 27072 9680 27084
rect 9732 27072 9738 27124
rect 11606 27072 11612 27124
rect 11664 27112 11670 27124
rect 11701 27115 11759 27121
rect 11701 27112 11713 27115
rect 11664 27084 11713 27112
rect 11664 27072 11670 27084
rect 11701 27081 11713 27084
rect 11747 27081 11759 27115
rect 11701 27075 11759 27081
rect 11882 27072 11888 27124
rect 11940 27112 11946 27124
rect 14458 27112 14464 27124
rect 11940 27084 14464 27112
rect 11940 27072 11946 27084
rect 14458 27072 14464 27084
rect 14516 27072 14522 27124
rect 14550 27072 14556 27124
rect 14608 27112 14614 27124
rect 18414 27112 18420 27124
rect 14608 27084 18420 27112
rect 14608 27072 14614 27084
rect 18414 27072 18420 27084
rect 18472 27072 18478 27124
rect 18690 27112 18696 27124
rect 18651 27084 18696 27112
rect 18690 27072 18696 27084
rect 18748 27072 18754 27124
rect 18877 27115 18935 27121
rect 18877 27081 18889 27115
rect 18923 27112 18935 27115
rect 18966 27112 18972 27124
rect 18923 27084 18972 27112
rect 18923 27081 18935 27084
rect 18877 27075 18935 27081
rect 18966 27072 18972 27084
rect 19024 27112 19030 27124
rect 20438 27112 20444 27124
rect 19024 27084 20444 27112
rect 19024 27072 19030 27084
rect 7374 27004 7380 27056
rect 7432 27004 7438 27056
rect 9858 27004 9864 27056
rect 9916 27004 9922 27056
rect 13538 27044 13544 27056
rect 13280 27016 13544 27044
rect 6178 26936 6184 26988
rect 6236 26976 6242 26988
rect 6457 26979 6515 26985
rect 6457 26976 6469 26979
rect 6236 26948 6469 26976
rect 6236 26936 6242 26948
rect 6457 26945 6469 26948
rect 6503 26945 6515 26979
rect 11882 26976 11888 26988
rect 11843 26948 11888 26976
rect 6457 26939 6515 26945
rect 11882 26936 11888 26948
rect 11940 26936 11946 26988
rect 6730 26908 6736 26920
rect 6691 26880 6736 26908
rect 6730 26868 6736 26880
rect 6788 26868 6794 26920
rect 8202 26908 8208 26920
rect 8115 26880 8208 26908
rect 8202 26868 8208 26880
rect 8260 26908 8266 26920
rect 9950 26908 9956 26920
rect 8260 26880 9956 26908
rect 8260 26868 8266 26880
rect 9950 26868 9956 26880
rect 10008 26868 10014 26920
rect 10318 26908 10324 26920
rect 10279 26880 10324 26908
rect 10318 26868 10324 26880
rect 10376 26868 10382 26920
rect 13280 26917 13308 27016
rect 13538 27004 13544 27016
rect 13596 27004 13602 27056
rect 14274 27004 14280 27056
rect 14332 27004 14338 27056
rect 14918 27004 14924 27056
rect 14976 27044 14982 27056
rect 18708 27044 18736 27072
rect 14976 27016 15976 27044
rect 14976 27004 14982 27016
rect 15654 26976 15660 26988
rect 15028 26948 15660 26976
rect 10597 26911 10655 26917
rect 10597 26877 10609 26911
rect 10643 26877 10655 26911
rect 13265 26911 13323 26917
rect 13265 26908 13277 26911
rect 10597 26871 10655 26877
rect 11624 26880 13277 26908
rect 9766 26732 9772 26784
rect 9824 26772 9830 26784
rect 10612 26772 10640 26871
rect 11624 26784 11652 26880
rect 13265 26877 13277 26880
rect 13311 26877 13323 26911
rect 13265 26871 13323 26877
rect 13541 26911 13599 26917
rect 13541 26877 13553 26911
rect 13587 26908 13599 26911
rect 14090 26908 14096 26920
rect 13587 26880 14096 26908
rect 13587 26877 13599 26880
rect 13541 26871 13599 26877
rect 14090 26868 14096 26880
rect 14148 26868 14154 26920
rect 15028 26917 15056 26948
rect 15654 26936 15660 26948
rect 15712 26936 15718 26988
rect 15948 26985 15976 27016
rect 16960 27016 18000 27044
rect 18708 27016 19748 27044
rect 16960 26988 16988 27016
rect 15841 26979 15899 26985
rect 15841 26945 15853 26979
rect 15887 26945 15899 26979
rect 15841 26939 15899 26945
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26945 15991 26979
rect 15933 26939 15991 26945
rect 15013 26911 15071 26917
rect 15013 26877 15025 26911
rect 15059 26877 15071 26911
rect 15856 26908 15884 26939
rect 16206 26936 16212 26988
rect 16264 26976 16270 26988
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16264 26948 16865 26976
rect 16264 26936 16270 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 16942 26936 16948 26988
rect 17000 26976 17006 26988
rect 17865 26979 17923 26985
rect 17000 26948 17045 26976
rect 17000 26936 17006 26948
rect 17865 26945 17877 26979
rect 17911 26945 17923 26979
rect 17972 26976 18000 27016
rect 18782 26976 18788 26988
rect 17972 26948 18788 26976
rect 17865 26939 17923 26945
rect 16574 26908 16580 26920
rect 15856 26880 16580 26908
rect 15013 26871 15071 26877
rect 16574 26868 16580 26880
rect 16632 26868 16638 26920
rect 17681 26911 17739 26917
rect 17681 26877 17693 26911
rect 17727 26877 17739 26911
rect 17880 26908 17908 26939
rect 18782 26936 18788 26948
rect 18840 26936 18846 26988
rect 19058 26976 19064 26988
rect 19019 26948 19064 26976
rect 19058 26936 19064 26948
rect 19116 26936 19122 26988
rect 19720 26985 19748 27016
rect 19904 26985 19932 27084
rect 20438 27072 20444 27084
rect 20496 27072 20502 27124
rect 21069 27115 21127 27121
rect 21069 27081 21081 27115
rect 21115 27112 21127 27115
rect 21174 27112 21180 27124
rect 21115 27084 21180 27112
rect 21115 27081 21127 27084
rect 21069 27075 21127 27081
rect 21174 27072 21180 27084
rect 21232 27112 21238 27124
rect 21818 27112 21824 27124
rect 21232 27084 21824 27112
rect 21232 27072 21238 27084
rect 21818 27072 21824 27084
rect 21876 27072 21882 27124
rect 27522 27072 27528 27124
rect 27580 27112 27586 27124
rect 28813 27115 28871 27121
rect 28813 27112 28825 27115
rect 27580 27084 28825 27112
rect 27580 27072 27586 27084
rect 28813 27081 28825 27084
rect 28859 27081 28871 27115
rect 28813 27075 28871 27081
rect 28902 27072 28908 27124
rect 28960 27112 28966 27124
rect 28960 27084 29868 27112
rect 28960 27072 28966 27084
rect 21266 27044 21272 27056
rect 21227 27016 21272 27044
rect 21266 27004 21272 27016
rect 21324 27004 21330 27056
rect 22738 27004 22744 27056
rect 22796 27004 22802 27056
rect 24397 27047 24455 27053
rect 24397 27013 24409 27047
rect 24443 27044 24455 27047
rect 24670 27044 24676 27056
rect 24443 27016 24676 27044
rect 24443 27013 24455 27016
rect 24397 27007 24455 27013
rect 24670 27004 24676 27016
rect 24728 27004 24734 27056
rect 24854 27004 24860 27056
rect 24912 27004 24918 27056
rect 29546 27044 29552 27056
rect 28566 27016 29552 27044
rect 29546 27004 29552 27016
rect 29604 27004 29610 27056
rect 29840 27053 29868 27084
rect 31294 27072 31300 27124
rect 31352 27112 31358 27124
rect 31573 27115 31631 27121
rect 31352 27084 31397 27112
rect 31352 27072 31358 27084
rect 31573 27081 31585 27115
rect 31619 27112 31631 27115
rect 32674 27112 32680 27124
rect 31619 27084 32680 27112
rect 31619 27081 31631 27084
rect 31573 27075 31631 27081
rect 32674 27072 32680 27084
rect 32732 27072 32738 27124
rect 32858 27072 32864 27124
rect 32916 27112 32922 27124
rect 32953 27115 33011 27121
rect 32953 27112 32965 27115
rect 32916 27084 32965 27112
rect 32916 27072 32922 27084
rect 32953 27081 32965 27084
rect 32999 27081 33011 27115
rect 32953 27075 33011 27081
rect 34701 27115 34759 27121
rect 34701 27081 34713 27115
rect 34747 27112 34759 27115
rect 34790 27112 34796 27124
rect 34747 27084 34796 27112
rect 34747 27081 34759 27084
rect 34701 27075 34759 27081
rect 34790 27072 34796 27084
rect 34848 27072 34854 27124
rect 37366 27112 37372 27124
rect 37327 27084 37372 27112
rect 37366 27072 37372 27084
rect 37424 27072 37430 27124
rect 29825 27047 29883 27053
rect 29825 27013 29837 27047
rect 29871 27013 29883 27047
rect 29825 27007 29883 27013
rect 29963 27047 30021 27053
rect 29963 27013 29975 27047
rect 30009 27044 30021 27047
rect 30374 27044 30380 27056
rect 30009 27016 30380 27044
rect 30009 27013 30021 27016
rect 29963 27007 30021 27013
rect 30374 27004 30380 27016
rect 30432 27004 30438 27056
rect 31389 27047 31447 27053
rect 31389 27044 31401 27047
rect 30484 27016 31401 27044
rect 19705 26979 19763 26985
rect 19705 26945 19717 26979
rect 19751 26945 19763 26979
rect 19705 26939 19763 26945
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26945 19947 26979
rect 19889 26939 19947 26945
rect 20806 26936 20812 26988
rect 20864 26976 20870 26988
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 20864 26948 21833 26976
rect 20864 26936 20870 26948
rect 21821 26945 21833 26948
rect 21867 26945 21879 26979
rect 29638 26976 29644 26988
rect 29599 26948 29644 26976
rect 21821 26939 21879 26945
rect 29638 26936 29644 26948
rect 29696 26936 29702 26988
rect 29730 26936 29736 26988
rect 29788 26976 29794 26988
rect 29788 26948 29833 26976
rect 29788 26936 29794 26948
rect 30190 26936 30196 26988
rect 30248 26976 30254 26988
rect 30484 26976 30512 27016
rect 31389 27013 31401 27016
rect 31435 27013 31447 27047
rect 31389 27007 31447 27013
rect 32398 27004 32404 27056
rect 32456 27044 32462 27056
rect 33965 27047 34023 27053
rect 33965 27044 33977 27047
rect 32456 27016 33977 27044
rect 32456 27004 32462 27016
rect 33965 27013 33977 27016
rect 34011 27013 34023 27047
rect 33965 27007 34023 27013
rect 34149 27047 34207 27053
rect 34149 27013 34161 27047
rect 34195 27044 34207 27047
rect 34330 27044 34336 27056
rect 34195 27016 34336 27044
rect 34195 27013 34207 27016
rect 34149 27007 34207 27013
rect 34330 27004 34336 27016
rect 34388 27044 34394 27056
rect 34514 27044 34520 27056
rect 34388 27016 34520 27044
rect 34388 27004 34394 27016
rect 34514 27004 34520 27016
rect 34572 27004 34578 27056
rect 30248 26948 30512 26976
rect 30248 26936 30254 26948
rect 31110 26936 31116 26988
rect 31168 26976 31174 26988
rect 31205 26979 31263 26985
rect 31205 26976 31217 26979
rect 31168 26948 31217 26976
rect 31168 26936 31174 26948
rect 31205 26945 31217 26948
rect 31251 26945 31263 26979
rect 31205 26939 31263 26945
rect 19521 26911 19579 26917
rect 19521 26908 19533 26911
rect 17880 26880 19533 26908
rect 17681 26871 17739 26877
rect 19521 26877 19533 26880
rect 19567 26877 19579 26911
rect 19794 26908 19800 26920
rect 19755 26880 19800 26908
rect 19521 26871 19579 26877
rect 17494 26840 17500 26852
rect 15304 26812 17500 26840
rect 11606 26772 11612 26784
rect 9824 26744 11612 26772
rect 9824 26732 9830 26744
rect 11606 26732 11612 26744
rect 11664 26732 11670 26784
rect 11698 26732 11704 26784
rect 11756 26772 11762 26784
rect 15304 26772 15332 26812
rect 17494 26800 17500 26812
rect 17552 26800 17558 26852
rect 17696 26840 17724 26871
rect 19794 26868 19800 26880
rect 19852 26868 19858 26920
rect 19981 26911 20039 26917
rect 19981 26877 19993 26911
rect 20027 26877 20039 26911
rect 19981 26871 20039 26877
rect 18874 26840 18880 26852
rect 17696 26812 18880 26840
rect 18874 26800 18880 26812
rect 18932 26800 18938 26852
rect 19058 26800 19064 26852
rect 19116 26840 19122 26852
rect 19996 26840 20024 26871
rect 22094 26868 22100 26920
rect 22152 26908 22158 26920
rect 24121 26911 24179 26917
rect 24121 26908 24133 26911
rect 22152 26880 22197 26908
rect 23216 26880 24133 26908
rect 22152 26868 22158 26880
rect 23216 26852 23244 26880
rect 24121 26877 24133 26880
rect 24167 26908 24179 26911
rect 25130 26908 25136 26920
rect 24167 26880 25136 26908
rect 24167 26877 24179 26880
rect 24121 26871 24179 26877
rect 25130 26868 25136 26880
rect 25188 26908 25194 26920
rect 27065 26911 27123 26917
rect 27065 26908 27077 26911
rect 25188 26880 27077 26908
rect 25188 26868 25194 26880
rect 27065 26877 27077 26880
rect 27111 26877 27123 26911
rect 27065 26871 27123 26877
rect 27341 26911 27399 26917
rect 27341 26877 27353 26911
rect 27387 26908 27399 26911
rect 27706 26908 27712 26920
rect 27387 26880 27712 26908
rect 27387 26877 27399 26880
rect 27341 26871 27399 26877
rect 27706 26868 27712 26880
rect 27764 26868 27770 26920
rect 30006 26868 30012 26920
rect 30064 26908 30070 26920
rect 30101 26911 30159 26917
rect 30101 26908 30113 26911
rect 30064 26880 30113 26908
rect 30064 26868 30070 26880
rect 30101 26877 30113 26880
rect 30147 26877 30159 26911
rect 30101 26871 30159 26877
rect 30282 26868 30288 26920
rect 30340 26908 30346 26920
rect 31220 26908 31248 26939
rect 31478 26936 31484 26988
rect 31536 26976 31542 26988
rect 32309 26979 32367 26985
rect 32309 26976 32321 26979
rect 31536 26948 32321 26976
rect 31536 26936 31542 26948
rect 32309 26945 32321 26948
rect 32355 26976 32367 26979
rect 32674 26976 32680 26988
rect 32355 26948 32680 26976
rect 32355 26945 32367 26948
rect 32309 26939 32367 26945
rect 32674 26936 32680 26948
rect 32732 26936 32738 26988
rect 33137 26979 33195 26985
rect 33137 26945 33149 26979
rect 33183 26945 33195 26979
rect 33410 26976 33416 26988
rect 33371 26948 33416 26976
rect 33137 26939 33195 26945
rect 31570 26908 31576 26920
rect 30340 26880 31576 26908
rect 30340 26868 30346 26880
rect 31570 26868 31576 26880
rect 31628 26868 31634 26920
rect 19116 26812 20024 26840
rect 19116 26800 19122 26812
rect 23198 26800 23204 26852
rect 23256 26800 23262 26852
rect 23566 26840 23572 26852
rect 23527 26812 23572 26840
rect 23566 26800 23572 26812
rect 23624 26800 23630 26852
rect 28350 26800 28356 26852
rect 28408 26840 28414 26852
rect 30834 26840 30840 26852
rect 28408 26812 30840 26840
rect 28408 26800 28414 26812
rect 30834 26800 30840 26812
rect 30892 26800 30898 26852
rect 31021 26843 31079 26849
rect 31021 26809 31033 26843
rect 31067 26840 31079 26843
rect 31202 26840 31208 26852
rect 31067 26812 31208 26840
rect 31067 26809 31079 26812
rect 31021 26803 31079 26809
rect 31202 26800 31208 26812
rect 31260 26840 31266 26852
rect 32490 26840 32496 26852
rect 31260 26812 32496 26840
rect 31260 26800 31266 26812
rect 32490 26800 32496 26812
rect 32548 26800 32554 26852
rect 33152 26840 33180 26939
rect 33410 26936 33416 26948
rect 33468 26936 33474 26988
rect 34609 26979 34667 26985
rect 34609 26945 34621 26979
rect 34655 26976 34667 26979
rect 34698 26976 34704 26988
rect 34655 26948 34704 26976
rect 34655 26945 34667 26948
rect 34609 26939 34667 26945
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 35253 26979 35311 26985
rect 35253 26945 35265 26979
rect 35299 26945 35311 26979
rect 35434 26976 35440 26988
rect 35395 26948 35440 26976
rect 35253 26939 35311 26945
rect 33226 26868 33232 26920
rect 33284 26908 33290 26920
rect 33321 26911 33379 26917
rect 33321 26908 33333 26911
rect 33284 26880 33333 26908
rect 33284 26868 33290 26880
rect 33321 26877 33333 26880
rect 33367 26908 33379 26911
rect 33778 26908 33784 26920
rect 33367 26880 33784 26908
rect 33367 26877 33379 26880
rect 33321 26871 33379 26877
rect 33778 26868 33784 26880
rect 33836 26868 33842 26920
rect 35268 26908 35296 26939
rect 35434 26936 35440 26948
rect 35492 26936 35498 26988
rect 37458 26976 37464 26988
rect 37419 26948 37464 26976
rect 37458 26936 37464 26948
rect 37516 26936 37522 26988
rect 35618 26908 35624 26920
rect 35268 26880 35624 26908
rect 35618 26868 35624 26880
rect 35676 26868 35682 26920
rect 33870 26840 33876 26852
rect 33152 26812 33876 26840
rect 33870 26800 33876 26812
rect 33928 26800 33934 26852
rect 15470 26772 15476 26784
rect 11756 26744 15332 26772
rect 15431 26744 15476 26772
rect 11756 26732 11762 26744
rect 15470 26732 15476 26744
rect 15528 26732 15534 26784
rect 15930 26732 15936 26784
rect 15988 26772 15994 26784
rect 16669 26775 16727 26781
rect 16669 26772 16681 26775
rect 15988 26744 16681 26772
rect 15988 26732 15994 26744
rect 16669 26741 16681 26744
rect 16715 26741 16727 26775
rect 18046 26772 18052 26784
rect 18007 26744 18052 26772
rect 16669 26735 16727 26741
rect 18046 26732 18052 26744
rect 18104 26732 18110 26784
rect 18322 26732 18328 26784
rect 18380 26772 18386 26784
rect 18509 26775 18567 26781
rect 18509 26772 18521 26775
rect 18380 26744 18521 26772
rect 18380 26732 18386 26744
rect 18509 26741 18521 26744
rect 18555 26741 18567 26775
rect 18509 26735 18567 26741
rect 18782 26732 18788 26784
rect 18840 26772 18846 26784
rect 20714 26772 20720 26784
rect 18840 26744 20720 26772
rect 18840 26732 18846 26744
rect 20714 26732 20720 26744
rect 20772 26732 20778 26784
rect 20898 26772 20904 26784
rect 20859 26744 20904 26772
rect 20898 26732 20904 26744
rect 20956 26732 20962 26784
rect 20990 26732 20996 26784
rect 21048 26772 21054 26784
rect 21085 26775 21143 26781
rect 21085 26772 21097 26775
rect 21048 26744 21097 26772
rect 21048 26732 21054 26744
rect 21085 26741 21097 26744
rect 21131 26741 21143 26775
rect 21085 26735 21143 26741
rect 25682 26732 25688 26784
rect 25740 26772 25746 26784
rect 25869 26775 25927 26781
rect 25869 26772 25881 26775
rect 25740 26744 25881 26772
rect 25740 26732 25746 26744
rect 25869 26741 25881 26744
rect 25915 26772 25927 26775
rect 28442 26772 28448 26784
rect 25915 26744 28448 26772
rect 25915 26741 25927 26744
rect 25869 26735 25927 26741
rect 28442 26732 28448 26744
rect 28500 26732 28506 26784
rect 29457 26775 29515 26781
rect 29457 26741 29469 26775
rect 29503 26772 29515 26775
rect 29822 26772 29828 26784
rect 29503 26744 29828 26772
rect 29503 26741 29515 26744
rect 29457 26735 29515 26741
rect 29822 26732 29828 26744
rect 29880 26732 29886 26784
rect 30650 26732 30656 26784
rect 30708 26772 30714 26784
rect 31478 26772 31484 26784
rect 30708 26744 31484 26772
rect 30708 26732 30714 26744
rect 31478 26732 31484 26744
rect 31536 26732 31542 26784
rect 32401 26775 32459 26781
rect 32401 26741 32413 26775
rect 32447 26772 32459 26775
rect 33318 26772 33324 26784
rect 32447 26744 33324 26772
rect 32447 26741 32459 26744
rect 32401 26735 32459 26741
rect 33318 26732 33324 26744
rect 33376 26732 33382 26784
rect 33413 26775 33471 26781
rect 33413 26741 33425 26775
rect 33459 26772 33471 26775
rect 34054 26772 34060 26784
rect 33459 26744 34060 26772
rect 33459 26741 33471 26744
rect 33413 26735 33471 26741
rect 34054 26732 34060 26744
rect 34112 26732 34118 26784
rect 34790 26732 34796 26784
rect 34848 26772 34854 26784
rect 35253 26775 35311 26781
rect 35253 26772 35265 26775
rect 34848 26744 35265 26772
rect 34848 26732 34854 26744
rect 35253 26741 35265 26744
rect 35299 26741 35311 26775
rect 35253 26735 35311 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 6730 26528 6736 26580
rect 6788 26568 6794 26580
rect 7009 26571 7067 26577
rect 7009 26568 7021 26571
rect 6788 26540 7021 26568
rect 6788 26528 6794 26540
rect 7009 26537 7021 26540
rect 7055 26537 7067 26571
rect 7009 26531 7067 26537
rect 10318 26528 10324 26580
rect 10376 26568 10382 26580
rect 10413 26571 10471 26577
rect 10413 26568 10425 26571
rect 10376 26540 10425 26568
rect 10376 26528 10382 26540
rect 10413 26537 10425 26540
rect 10459 26537 10471 26571
rect 10413 26531 10471 26537
rect 10870 26528 10876 26580
rect 10928 26568 10934 26580
rect 14550 26568 14556 26580
rect 10928 26540 14556 26568
rect 10928 26528 10934 26540
rect 14550 26528 14556 26540
rect 14608 26528 14614 26580
rect 15378 26568 15384 26580
rect 14752 26540 15384 26568
rect 7653 26503 7711 26509
rect 7653 26469 7665 26503
rect 7699 26469 7711 26503
rect 14752 26500 14780 26540
rect 15378 26528 15384 26540
rect 15436 26528 15442 26580
rect 18046 26528 18052 26580
rect 18104 26568 18110 26580
rect 18104 26540 21220 26568
rect 18104 26528 18110 26540
rect 15565 26503 15623 26509
rect 15565 26500 15577 26503
rect 7653 26463 7711 26469
rect 9968 26472 14780 26500
rect 14844 26472 15577 26500
rect 1854 26324 1860 26376
rect 1912 26364 1918 26376
rect 1949 26367 2007 26373
rect 1949 26364 1961 26367
rect 1912 26336 1961 26364
rect 1912 26324 1918 26336
rect 1949 26333 1961 26336
rect 1995 26333 2007 26367
rect 1949 26327 2007 26333
rect 7193 26367 7251 26373
rect 7193 26333 7205 26367
rect 7239 26364 7251 26367
rect 7668 26364 7696 26463
rect 8202 26432 8208 26444
rect 8163 26404 8208 26432
rect 8202 26392 8208 26404
rect 8260 26392 8266 26444
rect 8941 26435 8999 26441
rect 8941 26401 8953 26435
rect 8987 26432 8999 26435
rect 9861 26435 9919 26441
rect 9861 26432 9873 26435
rect 8987 26404 9873 26432
rect 8987 26401 8999 26404
rect 8941 26395 8999 26401
rect 9861 26401 9873 26404
rect 9907 26401 9919 26435
rect 9861 26395 9919 26401
rect 7239 26336 7696 26364
rect 8113 26367 8171 26373
rect 7239 26333 7251 26336
rect 7193 26327 7251 26333
rect 8113 26333 8125 26367
rect 8159 26364 8171 26367
rect 8956 26364 8984 26395
rect 9122 26364 9128 26376
rect 8159 26336 8984 26364
rect 9083 26336 9128 26364
rect 8159 26333 8171 26336
rect 8113 26327 8171 26333
rect 9122 26324 9128 26336
rect 9180 26324 9186 26376
rect 9306 26324 9312 26376
rect 9364 26364 9370 26376
rect 9968 26373 9996 26472
rect 14734 26432 14740 26444
rect 14695 26404 14740 26432
rect 14734 26392 14740 26404
rect 14792 26392 14798 26444
rect 9769 26367 9827 26373
rect 9769 26364 9781 26367
rect 9364 26336 9781 26364
rect 9364 26324 9370 26336
rect 9769 26333 9781 26336
rect 9815 26333 9827 26367
rect 9769 26327 9827 26333
rect 9953 26367 10011 26373
rect 9953 26333 9965 26367
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 10597 26367 10655 26373
rect 10597 26333 10609 26367
rect 10643 26333 10655 26367
rect 11974 26364 11980 26376
rect 11935 26336 11980 26364
rect 10597 26327 10655 26333
rect 8021 26299 8079 26305
rect 8021 26265 8033 26299
rect 8067 26296 8079 26299
rect 8938 26296 8944 26308
rect 8067 26268 8944 26296
rect 8067 26265 8079 26268
rect 8021 26259 8079 26265
rect 8938 26256 8944 26268
rect 8996 26256 9002 26308
rect 10612 26296 10640 26327
rect 11974 26324 11980 26336
rect 12032 26324 12038 26376
rect 12158 26364 12164 26376
rect 12119 26336 12164 26364
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 14093 26367 14151 26373
rect 14093 26333 14105 26367
rect 14139 26364 14151 26367
rect 14844 26364 14872 26472
rect 15565 26469 15577 26472
rect 15611 26469 15623 26503
rect 15565 26463 15623 26469
rect 16574 26460 16580 26512
rect 16632 26500 16638 26512
rect 16945 26503 17003 26509
rect 16945 26500 16957 26503
rect 16632 26472 16957 26500
rect 16632 26460 16638 26472
rect 16945 26469 16957 26472
rect 16991 26500 17003 26503
rect 16991 26472 18644 26500
rect 16991 26469 17003 26472
rect 16945 26463 17003 26469
rect 15470 26432 15476 26444
rect 14936 26404 15476 26432
rect 14936 26373 14964 26404
rect 15470 26392 15476 26404
rect 15528 26392 15534 26444
rect 16114 26432 16120 26444
rect 16075 26404 16120 26432
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 18506 26432 18512 26444
rect 18467 26404 18512 26432
rect 18506 26392 18512 26404
rect 18564 26392 18570 26444
rect 18616 26432 18644 26472
rect 19058 26460 19064 26512
rect 19116 26500 19122 26512
rect 19337 26503 19395 26509
rect 19337 26500 19349 26503
rect 19116 26472 19349 26500
rect 19116 26460 19122 26472
rect 19337 26469 19349 26472
rect 19383 26469 19395 26503
rect 19337 26463 19395 26469
rect 19794 26432 19800 26444
rect 18616 26404 19800 26432
rect 19794 26392 19800 26404
rect 19852 26392 19858 26444
rect 20806 26392 20812 26444
rect 20864 26432 20870 26444
rect 21085 26435 21143 26441
rect 21085 26432 21097 26435
rect 20864 26404 21097 26432
rect 20864 26392 20870 26404
rect 21085 26401 21097 26404
rect 21131 26401 21143 26435
rect 21085 26395 21143 26401
rect 14139 26336 14872 26364
rect 14921 26367 14979 26373
rect 14139 26333 14151 26336
rect 14093 26327 14151 26333
rect 14921 26333 14933 26367
rect 14967 26333 14979 26367
rect 14921 26327 14979 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26364 15163 26367
rect 15562 26364 15568 26376
rect 15151 26336 15568 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 15930 26364 15936 26376
rect 15891 26336 15936 26364
rect 15930 26324 15936 26336
rect 15988 26324 15994 26376
rect 16942 26324 16948 26376
rect 17000 26364 17006 26376
rect 17129 26367 17187 26373
rect 17129 26364 17141 26367
rect 17000 26336 17141 26364
rect 17000 26324 17006 26336
rect 17129 26333 17141 26336
rect 17175 26333 17187 26367
rect 18322 26364 18328 26376
rect 18283 26336 18328 26364
rect 17129 26327 17187 26333
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26364 18475 26367
rect 18874 26364 18880 26376
rect 18463 26336 18880 26364
rect 18463 26333 18475 26336
rect 18417 26327 18475 26333
rect 18874 26324 18880 26336
rect 18932 26324 18938 26376
rect 21192 26364 21220 26540
rect 21266 26528 21272 26580
rect 21324 26568 21330 26580
rect 24486 26568 24492 26580
rect 21324 26540 24492 26568
rect 21324 26528 21330 26540
rect 24486 26528 24492 26540
rect 24544 26568 24550 26580
rect 24765 26571 24823 26577
rect 24765 26568 24777 26571
rect 24544 26540 24777 26568
rect 24544 26528 24550 26540
rect 24765 26537 24777 26540
rect 24811 26537 24823 26571
rect 25866 26568 25872 26580
rect 25827 26540 25872 26568
rect 24765 26531 24823 26537
rect 25866 26528 25872 26540
rect 25924 26528 25930 26580
rect 26786 26568 26792 26580
rect 26747 26540 26792 26568
rect 26786 26528 26792 26540
rect 26844 26528 26850 26580
rect 31941 26571 31999 26577
rect 30024 26540 31754 26568
rect 22278 26500 22284 26512
rect 22239 26472 22284 26500
rect 22278 26460 22284 26472
rect 22336 26460 22342 26512
rect 26237 26503 26295 26509
rect 26237 26469 26249 26503
rect 26283 26500 26295 26503
rect 27798 26500 27804 26512
rect 26283 26472 27804 26500
rect 26283 26469 26295 26472
rect 26237 26463 26295 26469
rect 27798 26460 27804 26472
rect 27856 26460 27862 26512
rect 28261 26503 28319 26509
rect 28261 26469 28273 26503
rect 28307 26500 28319 26503
rect 28534 26500 28540 26512
rect 28307 26472 28540 26500
rect 28307 26469 28319 26472
rect 28261 26463 28319 26469
rect 28534 26460 28540 26472
rect 28592 26460 28598 26512
rect 25958 26432 25964 26444
rect 25919 26404 25964 26432
rect 25958 26392 25964 26404
rect 26016 26392 26022 26444
rect 27065 26435 27123 26441
rect 27065 26432 27077 26435
rect 26252 26404 27077 26432
rect 21729 26367 21787 26373
rect 21729 26364 21741 26367
rect 21192 26336 21741 26364
rect 21729 26333 21741 26336
rect 21775 26333 21787 26367
rect 21729 26327 21787 26333
rect 21818 26324 21824 26376
rect 21876 26364 21882 26376
rect 22554 26364 22560 26376
rect 21876 26336 22560 26364
rect 21876 26324 21882 26336
rect 22554 26324 22560 26336
rect 22612 26324 22618 26376
rect 22833 26367 22891 26373
rect 22833 26333 22845 26367
rect 22879 26333 22891 26367
rect 22833 26327 22891 26333
rect 23385 26367 23443 26373
rect 23385 26333 23397 26367
rect 23431 26333 23443 26367
rect 23385 26327 23443 26333
rect 23661 26367 23719 26373
rect 23661 26333 23673 26367
rect 23707 26364 23719 26367
rect 24118 26364 24124 26376
rect 23707 26336 24124 26364
rect 23707 26333 23719 26336
rect 23661 26327 23719 26333
rect 15470 26296 15476 26308
rect 9324 26268 10640 26296
rect 14292 26268 15476 26296
rect 9324 26237 9352 26268
rect 9309 26231 9367 26237
rect 9309 26197 9321 26231
rect 9355 26197 9367 26231
rect 12066 26228 12072 26240
rect 12027 26200 12072 26228
rect 9309 26191 9367 26197
rect 12066 26188 12072 26200
rect 12124 26188 12130 26240
rect 14292 26237 14320 26268
rect 15470 26256 15476 26268
rect 15528 26256 15534 26308
rect 15580 26296 15608 26324
rect 16025 26299 16083 26305
rect 16025 26296 16037 26299
rect 15580 26268 16037 26296
rect 16025 26265 16037 26268
rect 16071 26265 16083 26299
rect 16025 26259 16083 26265
rect 17788 26268 18092 26296
rect 14277 26231 14335 26237
rect 14277 26197 14289 26231
rect 14323 26197 14335 26231
rect 14277 26191 14335 26197
rect 15286 26188 15292 26240
rect 15344 26228 15350 26240
rect 17788 26228 17816 26268
rect 17954 26228 17960 26240
rect 15344 26200 17816 26228
rect 17915 26200 17960 26228
rect 15344 26188 15350 26200
rect 17954 26188 17960 26200
rect 18012 26188 18018 26240
rect 18064 26228 18092 26268
rect 20346 26256 20352 26308
rect 20404 26256 20410 26308
rect 20809 26299 20867 26305
rect 20809 26265 20821 26299
rect 20855 26296 20867 26299
rect 20855 26268 21588 26296
rect 20855 26265 20867 26268
rect 20809 26259 20867 26265
rect 21082 26228 21088 26240
rect 18064 26200 21088 26228
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 21560 26237 21588 26268
rect 22002 26256 22008 26308
rect 22060 26296 22066 26308
rect 22848 26296 22876 26327
rect 23400 26296 23428 26327
rect 24118 26324 24124 26336
rect 24176 26364 24182 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 24176 26336 24593 26364
rect 24176 26324 24182 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 24762 26324 24768 26376
rect 24820 26364 24826 26376
rect 25777 26367 25835 26373
rect 25777 26364 25789 26367
rect 24820 26336 25789 26364
rect 24820 26324 24826 26336
rect 25777 26333 25789 26336
rect 25823 26333 25835 26367
rect 26050 26364 26056 26376
rect 26011 26336 26056 26364
rect 25777 26327 25835 26333
rect 26050 26324 26056 26336
rect 26108 26324 26114 26376
rect 23474 26296 23480 26308
rect 22060 26268 22876 26296
rect 23387 26268 23480 26296
rect 22060 26256 22066 26268
rect 23474 26256 23480 26268
rect 23532 26296 23538 26308
rect 24394 26296 24400 26308
rect 23532 26268 24400 26296
rect 23532 26256 23538 26268
rect 24394 26256 24400 26268
rect 24452 26256 24458 26308
rect 21545 26231 21603 26237
rect 21545 26197 21557 26231
rect 21591 26197 21603 26231
rect 21545 26191 21603 26197
rect 25958 26188 25964 26240
rect 26016 26228 26022 26240
rect 26252 26228 26280 26404
rect 27065 26401 27077 26404
rect 27111 26401 27123 26435
rect 27065 26395 27123 26401
rect 27249 26435 27307 26441
rect 27249 26401 27261 26435
rect 27295 26432 27307 26435
rect 28442 26432 28448 26444
rect 27295 26404 28448 26432
rect 27295 26401 27307 26404
rect 27249 26395 27307 26401
rect 28442 26392 28448 26404
rect 28500 26392 28506 26444
rect 28718 26432 28724 26444
rect 28679 26404 28724 26432
rect 28718 26392 28724 26404
rect 28776 26392 28782 26444
rect 28905 26435 28963 26441
rect 28905 26401 28917 26435
rect 28951 26432 28963 26435
rect 29914 26432 29920 26444
rect 28951 26404 29920 26432
rect 28951 26401 28963 26404
rect 28905 26395 28963 26401
rect 29914 26392 29920 26404
rect 29972 26392 29978 26444
rect 26418 26324 26424 26376
rect 26476 26364 26482 26376
rect 26973 26367 27031 26373
rect 26973 26364 26985 26367
rect 26476 26336 26985 26364
rect 26476 26324 26482 26336
rect 26973 26333 26985 26336
rect 27019 26333 27031 26367
rect 26973 26327 27031 26333
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 26326 26256 26332 26308
rect 26384 26296 26390 26308
rect 27172 26296 27200 26327
rect 27982 26324 27988 26376
rect 28040 26364 28046 26376
rect 28629 26367 28687 26373
rect 28629 26364 28641 26367
rect 28040 26336 28641 26364
rect 28040 26324 28046 26336
rect 28629 26333 28641 26336
rect 28675 26333 28687 26367
rect 28629 26327 28687 26333
rect 27522 26296 27528 26308
rect 26384 26268 27528 26296
rect 26384 26256 26390 26268
rect 27522 26256 27528 26268
rect 27580 26296 27586 26308
rect 27890 26296 27896 26308
rect 27580 26268 27896 26296
rect 27580 26256 27586 26268
rect 27890 26256 27896 26268
rect 27948 26256 27954 26308
rect 28902 26256 28908 26308
rect 28960 26296 28966 26308
rect 30024 26296 30052 26540
rect 30834 26460 30840 26512
rect 30892 26500 30898 26512
rect 31205 26503 31263 26509
rect 31205 26500 31217 26503
rect 30892 26472 31217 26500
rect 30892 26460 30898 26472
rect 31205 26469 31217 26472
rect 31251 26469 31263 26503
rect 31726 26500 31754 26540
rect 31941 26537 31953 26571
rect 31987 26568 31999 26571
rect 32398 26568 32404 26580
rect 31987 26540 32404 26568
rect 31987 26537 31999 26540
rect 31941 26531 31999 26537
rect 32398 26528 32404 26540
rect 32456 26528 32462 26580
rect 34422 26528 34428 26580
rect 34480 26568 34486 26580
rect 34701 26571 34759 26577
rect 34701 26568 34713 26571
rect 34480 26540 34713 26568
rect 34480 26528 34486 26540
rect 34701 26537 34713 26540
rect 34747 26537 34759 26571
rect 34701 26531 34759 26537
rect 34149 26503 34207 26509
rect 31726 26472 32352 26500
rect 31205 26463 31263 26469
rect 30098 26392 30104 26444
rect 30156 26432 30162 26444
rect 30156 26404 30201 26432
rect 30156 26392 30162 26404
rect 30282 26373 30288 26376
rect 30259 26367 30288 26373
rect 30259 26333 30271 26367
rect 30259 26327 30288 26333
rect 30282 26324 30288 26327
rect 30340 26324 30346 26376
rect 30558 26324 30564 26376
rect 30616 26364 30622 26376
rect 31389 26367 31447 26373
rect 30616 26336 30660 26364
rect 30616 26324 30622 26336
rect 31389 26333 31401 26367
rect 31435 26364 31447 26367
rect 31478 26364 31484 26376
rect 31435 26336 31484 26364
rect 31435 26333 31447 26336
rect 31389 26327 31447 26333
rect 31478 26324 31484 26336
rect 31536 26324 31542 26376
rect 32122 26364 32128 26376
rect 32083 26336 32128 26364
rect 32122 26324 32128 26336
rect 32180 26324 32186 26376
rect 32324 26373 32352 26472
rect 34149 26469 34161 26503
rect 34195 26500 34207 26503
rect 34606 26500 34612 26512
rect 34195 26472 34612 26500
rect 34195 26469 34207 26472
rect 34149 26463 34207 26469
rect 34606 26460 34612 26472
rect 34664 26460 34670 26512
rect 32585 26435 32643 26441
rect 32585 26401 32597 26435
rect 32631 26432 32643 26435
rect 33318 26432 33324 26444
rect 32631 26404 33324 26432
rect 32631 26401 32643 26404
rect 32585 26395 32643 26401
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 34790 26432 34796 26444
rect 33796 26404 34796 26432
rect 32309 26367 32367 26373
rect 32309 26333 32321 26367
rect 32355 26333 32367 26367
rect 32309 26327 32367 26333
rect 33597 26367 33655 26373
rect 33597 26333 33609 26367
rect 33643 26364 33655 26367
rect 33686 26364 33692 26376
rect 33643 26336 33692 26364
rect 33643 26333 33655 26336
rect 33597 26327 33655 26333
rect 33686 26324 33692 26336
rect 33744 26324 33750 26376
rect 33796 26373 33824 26404
rect 34790 26392 34796 26404
rect 34848 26392 34854 26444
rect 34900 26404 35756 26432
rect 33781 26367 33839 26373
rect 33781 26333 33793 26367
rect 33827 26333 33839 26367
rect 33962 26364 33968 26376
rect 33923 26336 33968 26364
rect 33781 26327 33839 26333
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34054 26324 34060 26376
rect 34112 26364 34118 26376
rect 34900 26373 34928 26404
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34112 26336 34897 26364
rect 34112 26324 34118 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 34977 26367 35035 26373
rect 34977 26333 34989 26367
rect 35023 26364 35035 26367
rect 35434 26364 35440 26376
rect 35023 26336 35440 26364
rect 35023 26333 35035 26336
rect 34977 26327 35035 26333
rect 30377 26299 30435 26305
rect 30377 26296 30389 26299
rect 28960 26268 30389 26296
rect 28960 26256 28966 26268
rect 30377 26265 30389 26268
rect 30423 26265 30435 26299
rect 30377 26259 30435 26265
rect 30466 26256 30472 26308
rect 30524 26296 30530 26308
rect 32214 26296 32220 26308
rect 30524 26268 30569 26296
rect 32175 26268 32220 26296
rect 30524 26256 30530 26268
rect 32214 26256 32220 26268
rect 32272 26256 32278 26308
rect 32490 26305 32496 26308
rect 32447 26299 32496 26305
rect 32447 26296 32459 26299
rect 32403 26268 32459 26296
rect 32447 26265 32459 26268
rect 32493 26265 32496 26299
rect 32447 26259 32496 26265
rect 32490 26256 32496 26259
rect 32548 26296 32554 26308
rect 33226 26296 33232 26308
rect 32548 26268 33232 26296
rect 32548 26256 32554 26268
rect 33226 26256 33232 26268
rect 33284 26256 33290 26308
rect 33870 26296 33876 26308
rect 33831 26268 33876 26296
rect 33870 26256 33876 26268
rect 33928 26296 33934 26308
rect 34992 26296 35020 26327
rect 35434 26324 35440 26336
rect 35492 26324 35498 26376
rect 35526 26324 35532 26376
rect 35584 26364 35590 26376
rect 35728 26373 35756 26404
rect 35713 26367 35771 26373
rect 35584 26336 35629 26364
rect 35584 26324 35590 26336
rect 35713 26333 35725 26367
rect 35759 26364 35771 26367
rect 35802 26364 35808 26376
rect 35759 26336 35808 26364
rect 35759 26333 35771 26336
rect 35713 26327 35771 26333
rect 35802 26324 35808 26336
rect 35860 26324 35866 26376
rect 36262 26324 36268 26376
rect 36320 26364 36326 26376
rect 37001 26367 37059 26373
rect 37001 26364 37013 26367
rect 36320 26336 37013 26364
rect 36320 26324 36326 26336
rect 37001 26333 37013 26336
rect 37047 26333 37059 26367
rect 37001 26327 37059 26333
rect 37829 26367 37887 26373
rect 37829 26333 37841 26367
rect 37875 26364 37887 26367
rect 37918 26364 37924 26376
rect 37875 26336 37924 26364
rect 37875 26333 37887 26336
rect 37829 26327 37887 26333
rect 37918 26324 37924 26336
rect 37976 26324 37982 26376
rect 35618 26296 35624 26308
rect 33928 26268 35020 26296
rect 35579 26268 35624 26296
rect 33928 26256 33934 26268
rect 35618 26256 35624 26268
rect 35676 26256 35682 26308
rect 26016 26200 26280 26228
rect 26016 26188 26022 26200
rect 30558 26188 30564 26240
rect 30616 26228 30622 26240
rect 30745 26231 30803 26237
rect 30745 26228 30757 26231
rect 30616 26200 30757 26228
rect 30616 26188 30622 26200
rect 30745 26197 30757 26200
rect 30791 26197 30803 26231
rect 30745 26191 30803 26197
rect 30834 26188 30840 26240
rect 30892 26228 30898 26240
rect 37274 26228 37280 26240
rect 30892 26200 37280 26228
rect 30892 26188 30898 26200
rect 37274 26188 37280 26200
rect 37332 26188 37338 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 7374 26024 7380 26036
rect 7335 25996 7380 26024
rect 7374 25984 7380 25996
rect 7432 25984 7438 26036
rect 9858 25984 9864 26036
rect 9916 26024 9922 26036
rect 10137 26027 10195 26033
rect 10137 26024 10149 26027
rect 9916 25996 10149 26024
rect 9916 25984 9922 25996
rect 10137 25993 10149 25996
rect 10183 25993 10195 26027
rect 14274 26024 14280 26036
rect 14235 25996 14280 26024
rect 10137 25987 10195 25993
rect 14274 25984 14280 25996
rect 14332 25984 14338 26036
rect 15562 26024 15568 26036
rect 15523 25996 15568 26024
rect 15562 25984 15568 25996
rect 15620 25984 15626 26036
rect 18322 26024 18328 26036
rect 16500 25996 18328 26024
rect 9401 25959 9459 25965
rect 9401 25925 9413 25959
rect 9447 25956 9459 25959
rect 11790 25956 11796 25968
rect 9447 25928 11796 25956
rect 9447 25925 9459 25928
rect 9401 25919 9459 25925
rect 11790 25916 11796 25928
rect 11848 25916 11854 25968
rect 11968 25959 12026 25965
rect 11968 25925 11980 25959
rect 12014 25956 12026 25959
rect 12066 25956 12072 25968
rect 12014 25928 12072 25956
rect 12014 25925 12026 25928
rect 11968 25919 12026 25925
rect 12066 25916 12072 25928
rect 12124 25916 12130 25968
rect 15286 25956 15292 25968
rect 12406 25928 15292 25956
rect 1854 25888 1860 25900
rect 1815 25860 1860 25888
rect 1854 25848 1860 25860
rect 1912 25848 1918 25900
rect 7282 25888 7288 25900
rect 7243 25860 7288 25888
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 9122 25848 9128 25900
rect 9180 25888 9186 25900
rect 9309 25891 9367 25897
rect 9309 25888 9321 25891
rect 9180 25860 9321 25888
rect 9180 25848 9186 25860
rect 9309 25857 9321 25860
rect 9355 25857 9367 25891
rect 9309 25851 9367 25857
rect 9585 25891 9643 25897
rect 9585 25857 9597 25891
rect 9631 25888 9643 25891
rect 10134 25888 10140 25900
rect 9631 25860 10140 25888
rect 9631 25857 9643 25860
rect 9585 25851 9643 25857
rect 10134 25848 10140 25860
rect 10192 25848 10198 25900
rect 10226 25848 10232 25900
rect 10284 25888 10290 25900
rect 10284 25860 10329 25888
rect 10284 25848 10290 25860
rect 11606 25848 11612 25900
rect 11664 25888 11670 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 11664 25860 11713 25888
rect 11664 25848 11670 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 12406 25888 12434 25928
rect 15286 25916 15292 25928
rect 15344 25916 15350 25968
rect 15470 25916 15476 25968
rect 15528 25956 15534 25968
rect 16390 25956 16396 25968
rect 15528 25928 16396 25956
rect 15528 25916 15534 25928
rect 16390 25916 16396 25928
rect 16448 25916 16454 25968
rect 11701 25851 11759 25857
rect 11808 25860 12434 25888
rect 14185 25891 14243 25897
rect 2041 25823 2099 25829
rect 2041 25789 2053 25823
rect 2087 25820 2099 25823
rect 2774 25820 2780 25832
rect 2087 25792 2780 25820
rect 2087 25789 2099 25792
rect 2041 25783 2099 25789
rect 2774 25780 2780 25792
rect 2832 25780 2838 25832
rect 2866 25780 2872 25832
rect 2924 25820 2930 25832
rect 2924 25792 2969 25820
rect 2924 25780 2930 25792
rect 6546 25780 6552 25832
rect 6604 25820 6610 25832
rect 11808 25820 11836 25860
rect 14185 25857 14197 25891
rect 14231 25888 14243 25891
rect 14826 25888 14832 25900
rect 14231 25860 14832 25888
rect 14231 25857 14243 25860
rect 14185 25851 14243 25857
rect 14826 25848 14832 25860
rect 14884 25848 14890 25900
rect 15102 25888 15108 25900
rect 15063 25860 15108 25888
rect 15102 25848 15108 25860
rect 15160 25848 15166 25900
rect 15838 25888 15844 25900
rect 15751 25860 15844 25888
rect 15838 25848 15844 25860
rect 15896 25888 15902 25900
rect 16500 25888 16528 25996
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 18417 26027 18475 26033
rect 18417 25993 18429 26027
rect 18463 26024 18475 26027
rect 18598 26024 18604 26036
rect 18463 25996 18604 26024
rect 18463 25993 18475 25996
rect 18417 25987 18475 25993
rect 18598 25984 18604 25996
rect 18656 25984 18662 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 22465 26027 22523 26033
rect 22152 25996 22197 26024
rect 22152 25984 22158 25996
rect 22465 25993 22477 26027
rect 22511 26024 22523 26027
rect 23566 26024 23572 26036
rect 22511 25996 23572 26024
rect 22511 25993 22523 25996
rect 22465 25987 22523 25993
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 24854 26024 24860 26036
rect 24815 25996 24860 26024
rect 24854 25984 24860 25996
rect 24912 25984 24918 26036
rect 27341 26027 27399 26033
rect 27341 26024 27353 26027
rect 26436 25996 27353 26024
rect 26436 25968 26464 25996
rect 27341 25993 27353 25996
rect 27387 25993 27399 26027
rect 27890 26024 27896 26036
rect 27851 25996 27896 26024
rect 27341 25987 27399 25993
rect 16574 25916 16580 25968
rect 16632 25956 16638 25968
rect 16945 25959 17003 25965
rect 16945 25956 16957 25959
rect 16632 25928 16957 25956
rect 16632 25916 16638 25928
rect 16945 25925 16957 25928
rect 16991 25925 17003 25959
rect 16945 25919 17003 25925
rect 17402 25916 17408 25968
rect 17460 25916 17466 25968
rect 20898 25956 20904 25968
rect 18248 25928 20904 25956
rect 16666 25888 16672 25900
rect 15896 25860 16528 25888
rect 16627 25860 16672 25888
rect 15896 25848 15902 25860
rect 16666 25848 16672 25860
rect 16724 25848 16730 25900
rect 6604 25792 11836 25820
rect 6604 25780 6610 25792
rect 15378 25780 15384 25832
rect 15436 25820 15442 25832
rect 15565 25823 15623 25829
rect 15565 25820 15577 25823
rect 15436 25792 15577 25820
rect 15436 25780 15442 25792
rect 15565 25789 15577 25792
rect 15611 25789 15623 25823
rect 15565 25783 15623 25789
rect 15749 25823 15807 25829
rect 15749 25789 15761 25823
rect 15795 25820 15807 25823
rect 16206 25820 16212 25832
rect 15795 25792 16212 25820
rect 15795 25789 15807 25792
rect 15749 25783 15807 25789
rect 15580 25752 15608 25783
rect 16206 25780 16212 25792
rect 16264 25780 16270 25832
rect 18248 25820 18276 25928
rect 20898 25916 20904 25928
rect 20956 25916 20962 25968
rect 21069 25959 21127 25965
rect 21069 25925 21081 25959
rect 21115 25956 21127 25959
rect 21115 25928 21220 25956
rect 21115 25925 21127 25928
rect 21069 25919 21127 25925
rect 19429 25891 19487 25897
rect 19429 25857 19441 25891
rect 19475 25888 19487 25891
rect 20254 25888 20260 25900
rect 19475 25860 20260 25888
rect 19475 25857 19487 25860
rect 19429 25851 19487 25857
rect 20254 25848 20260 25860
rect 20312 25848 20318 25900
rect 20441 25891 20499 25897
rect 20441 25857 20453 25891
rect 20487 25857 20499 25891
rect 21192 25888 21220 25928
rect 21266 25916 21272 25968
rect 21324 25956 21330 25968
rect 26418 25956 26424 25968
rect 21324 25928 21369 25956
rect 23216 25928 25636 25956
rect 26379 25928 26424 25956
rect 21324 25916 21330 25928
rect 22278 25888 22284 25900
rect 21192 25860 22284 25888
rect 20441 25851 20499 25857
rect 16316 25792 18276 25820
rect 20456 25820 20484 25851
rect 22278 25848 22284 25860
rect 22336 25848 22342 25900
rect 22557 25891 22615 25897
rect 22557 25857 22569 25891
rect 22603 25888 22615 25891
rect 23109 25891 23167 25897
rect 23109 25888 23121 25891
rect 22603 25860 23121 25888
rect 22603 25857 22615 25860
rect 22557 25851 22615 25857
rect 23109 25857 23121 25860
rect 23155 25857 23167 25891
rect 23109 25851 23167 25857
rect 22738 25820 22744 25832
rect 20456 25792 22744 25820
rect 16316 25752 16344 25792
rect 22738 25780 22744 25792
rect 22796 25780 22802 25832
rect 15580 25724 16344 25752
rect 19613 25755 19671 25761
rect 19613 25721 19625 25755
rect 19659 25752 19671 25755
rect 20714 25752 20720 25764
rect 19659 25724 20720 25752
rect 19659 25721 19671 25724
rect 19613 25715 19671 25721
rect 20714 25712 20720 25724
rect 20772 25712 20778 25764
rect 20806 25712 20812 25764
rect 20864 25752 20870 25764
rect 20901 25755 20959 25761
rect 20901 25752 20913 25755
rect 20864 25724 20913 25752
rect 20864 25712 20870 25724
rect 20901 25721 20913 25724
rect 20947 25721 20959 25755
rect 20901 25715 20959 25721
rect 21450 25712 21456 25764
rect 21508 25752 21514 25764
rect 23216 25752 23244 25928
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25888 23351 25891
rect 23477 25891 23535 25897
rect 23339 25860 23428 25888
rect 23339 25857 23351 25860
rect 23293 25851 23351 25857
rect 21508 25724 23244 25752
rect 23400 25752 23428 25860
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 23492 25820 23520 25851
rect 23566 25848 23572 25900
rect 23624 25888 23630 25900
rect 24118 25888 24124 25900
rect 23624 25860 23669 25888
rect 24079 25860 24124 25888
rect 23624 25848 23630 25860
rect 24118 25848 24124 25860
rect 24176 25848 24182 25900
rect 24578 25848 24584 25900
rect 24636 25888 24642 25900
rect 24765 25891 24823 25897
rect 24765 25888 24777 25891
rect 24636 25860 24777 25888
rect 24636 25848 24642 25860
rect 24765 25857 24777 25860
rect 24811 25857 24823 25891
rect 24765 25851 24823 25857
rect 25409 25891 25467 25897
rect 25409 25857 25421 25891
rect 25455 25888 25467 25891
rect 25498 25888 25504 25900
rect 25455 25860 25504 25888
rect 25455 25857 25467 25860
rect 25409 25851 25467 25857
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 25608 25897 25636 25928
rect 26418 25916 26424 25928
rect 26476 25916 26482 25968
rect 26973 25959 27031 25965
rect 26973 25925 26985 25959
rect 27019 25925 27031 25959
rect 26973 25919 27031 25925
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25888 26295 25891
rect 26326 25888 26332 25900
rect 26283 25860 26332 25888
rect 26283 25857 26295 25860
rect 26237 25851 26295 25857
rect 26326 25848 26332 25860
rect 26384 25848 26390 25900
rect 25958 25820 25964 25832
rect 23492 25792 25964 25820
rect 25958 25780 25964 25792
rect 26016 25780 26022 25832
rect 26142 25780 26148 25832
rect 26200 25820 26206 25832
rect 26988 25820 27016 25919
rect 27062 25916 27068 25968
rect 27120 25956 27126 25968
rect 27173 25959 27231 25965
rect 27173 25956 27185 25959
rect 27120 25928 27185 25956
rect 27120 25916 27126 25928
rect 27173 25925 27185 25928
rect 27219 25925 27231 25959
rect 27173 25919 27231 25925
rect 27356 25888 27384 25987
rect 27890 25984 27896 25996
rect 27948 25984 27954 26036
rect 30926 26024 30932 26036
rect 28092 25996 30932 26024
rect 28092 25965 28120 25996
rect 30926 25984 30932 25996
rect 30984 25984 30990 26036
rect 31202 25984 31208 26036
rect 31260 26024 31266 26036
rect 32030 26024 32036 26036
rect 31260 25996 32036 26024
rect 31260 25984 31266 25996
rect 32030 25984 32036 25996
rect 32088 25984 32094 26036
rect 33413 26027 33471 26033
rect 33413 25993 33425 26027
rect 33459 26024 33471 26027
rect 33594 26024 33600 26036
rect 33459 25996 33600 26024
rect 33459 25993 33471 25996
rect 33413 25987 33471 25993
rect 33594 25984 33600 25996
rect 33652 26024 33658 26036
rect 33962 26024 33968 26036
rect 33652 25996 33968 26024
rect 33652 25984 33658 25996
rect 33962 25984 33968 25996
rect 34020 25984 34026 26036
rect 35434 25984 35440 26036
rect 35492 26024 35498 26036
rect 36081 26027 36139 26033
rect 36081 26024 36093 26027
rect 35492 25996 36093 26024
rect 35492 25984 35498 25996
rect 36081 25993 36093 25996
rect 36127 25993 36139 26027
rect 36081 25987 36139 25993
rect 28077 25959 28135 25965
rect 28077 25925 28089 25959
rect 28123 25925 28135 25959
rect 30742 25956 30748 25968
rect 28077 25919 28135 25925
rect 29932 25928 30748 25956
rect 29932 25900 29960 25928
rect 30742 25916 30748 25928
rect 30800 25916 30806 25968
rect 31386 25916 31392 25968
rect 31444 25956 31450 25968
rect 33781 25959 33839 25965
rect 33781 25956 33793 25959
rect 31444 25928 33793 25956
rect 31444 25916 31450 25928
rect 33781 25925 33793 25928
rect 33827 25925 33839 25959
rect 34606 25956 34612 25968
rect 34567 25928 34612 25956
rect 33781 25919 33839 25925
rect 34606 25916 34612 25928
rect 34664 25916 34670 25968
rect 35342 25916 35348 25968
rect 35400 25916 35406 25968
rect 27801 25891 27859 25897
rect 27801 25888 27813 25891
rect 27356 25860 27813 25888
rect 27801 25857 27813 25860
rect 27847 25857 27859 25891
rect 28810 25888 28816 25900
rect 28771 25860 28816 25888
rect 27801 25851 27859 25857
rect 28810 25848 28816 25860
rect 28868 25848 28874 25900
rect 29914 25888 29920 25900
rect 29827 25860 29920 25888
rect 29914 25848 29920 25860
rect 29972 25848 29978 25900
rect 30190 25888 30196 25900
rect 30151 25860 30196 25888
rect 30190 25848 30196 25860
rect 30248 25848 30254 25900
rect 30650 25888 30656 25900
rect 30563 25860 30656 25888
rect 30650 25848 30656 25860
rect 30708 25888 30714 25900
rect 31294 25888 31300 25900
rect 30708 25860 31300 25888
rect 30708 25848 30714 25860
rect 31294 25848 31300 25860
rect 31352 25848 31358 25900
rect 31570 25848 31576 25900
rect 31628 25888 31634 25900
rect 32401 25891 32459 25897
rect 32401 25888 32413 25891
rect 31628 25860 32413 25888
rect 31628 25848 31634 25860
rect 32401 25857 32413 25860
rect 32447 25857 32459 25891
rect 32401 25851 32459 25857
rect 32674 25848 32680 25900
rect 32732 25888 32738 25900
rect 33597 25891 33655 25897
rect 33597 25888 33609 25891
rect 32732 25860 33609 25888
rect 32732 25848 32738 25860
rect 33597 25857 33609 25860
rect 33643 25857 33655 25891
rect 33597 25851 33655 25857
rect 33873 25891 33931 25897
rect 33873 25857 33885 25891
rect 33919 25857 33931 25891
rect 34330 25888 34336 25900
rect 34291 25860 34336 25888
rect 33873 25851 33931 25857
rect 28629 25823 28687 25829
rect 28629 25820 28641 25823
rect 26200 25792 27016 25820
rect 27908 25792 28641 25820
rect 26200 25780 26206 25792
rect 23474 25752 23480 25764
rect 23400 25724 23480 25752
rect 21508 25712 21514 25724
rect 23474 25712 23480 25724
rect 23532 25712 23538 25764
rect 24305 25755 24363 25761
rect 24305 25721 24317 25755
rect 24351 25752 24363 25755
rect 25590 25752 25596 25764
rect 24351 25724 25596 25752
rect 24351 25721 24363 25724
rect 24305 25715 24363 25721
rect 25590 25712 25596 25724
rect 25648 25712 25654 25764
rect 25976 25752 26004 25780
rect 27908 25752 27936 25792
rect 28629 25789 28641 25792
rect 28675 25820 28687 25823
rect 28902 25820 28908 25832
rect 28675 25792 28908 25820
rect 28675 25789 28687 25792
rect 28629 25783 28687 25789
rect 28902 25780 28908 25792
rect 28960 25780 28966 25832
rect 30006 25780 30012 25832
rect 30064 25820 30070 25832
rect 30374 25820 30380 25832
rect 30064 25792 30380 25820
rect 30064 25780 30070 25792
rect 30374 25780 30380 25792
rect 30432 25820 30438 25832
rect 30926 25820 30932 25832
rect 30432 25792 30932 25820
rect 30432 25780 30438 25792
rect 30926 25780 30932 25792
rect 30984 25780 30990 25832
rect 32030 25780 32036 25832
rect 32088 25820 32094 25832
rect 32125 25823 32183 25829
rect 32125 25820 32137 25823
rect 32088 25792 32137 25820
rect 32088 25780 32094 25792
rect 32125 25789 32137 25792
rect 32171 25820 32183 25823
rect 33410 25820 33416 25832
rect 32171 25792 33416 25820
rect 32171 25789 32183 25792
rect 32125 25783 32183 25789
rect 33410 25780 33416 25792
rect 33468 25780 33474 25832
rect 33888 25820 33916 25851
rect 34330 25848 34336 25860
rect 34388 25848 34394 25900
rect 37274 25888 37280 25900
rect 37235 25860 37280 25888
rect 37274 25848 37280 25860
rect 37332 25888 37338 25900
rect 37642 25888 37648 25900
rect 37332 25860 37648 25888
rect 37332 25848 37338 25860
rect 37642 25848 37648 25860
rect 37700 25848 37706 25900
rect 35618 25820 35624 25832
rect 33888 25792 35624 25820
rect 35618 25780 35624 25792
rect 35676 25780 35682 25832
rect 28074 25752 28080 25764
rect 25976 25724 27936 25752
rect 28035 25724 28080 25752
rect 28074 25712 28080 25724
rect 28132 25712 28138 25764
rect 9585 25687 9643 25693
rect 9585 25653 9597 25687
rect 9631 25684 9643 25687
rect 9674 25684 9680 25696
rect 9631 25656 9680 25684
rect 9631 25653 9643 25656
rect 9585 25647 9643 25653
rect 9674 25644 9680 25656
rect 9732 25644 9738 25696
rect 13078 25684 13084 25696
rect 13039 25656 13084 25684
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 15013 25687 15071 25693
rect 15013 25653 15025 25687
rect 15059 25684 15071 25687
rect 18230 25684 18236 25696
rect 15059 25656 18236 25684
rect 15059 25653 15071 25656
rect 15013 25647 15071 25653
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 20254 25684 20260 25696
rect 19484 25656 20260 25684
rect 19484 25644 19490 25656
rect 20254 25644 20260 25656
rect 20312 25644 20318 25696
rect 20990 25644 20996 25696
rect 21048 25684 21054 25696
rect 21085 25687 21143 25693
rect 21085 25684 21097 25687
rect 21048 25656 21097 25684
rect 21048 25644 21054 25656
rect 21085 25653 21097 25656
rect 21131 25684 21143 25687
rect 22002 25684 22008 25696
rect 21131 25656 22008 25684
rect 21131 25653 21143 25656
rect 21085 25647 21143 25653
rect 22002 25644 22008 25656
rect 22060 25644 22066 25696
rect 25406 25644 25412 25696
rect 25464 25684 25470 25696
rect 25501 25687 25559 25693
rect 25501 25684 25513 25687
rect 25464 25656 25513 25684
rect 25464 25644 25470 25656
rect 25501 25653 25513 25656
rect 25547 25653 25559 25687
rect 25501 25647 25559 25653
rect 26053 25687 26111 25693
rect 26053 25653 26065 25687
rect 26099 25684 26111 25687
rect 26970 25684 26976 25696
rect 26099 25656 26976 25684
rect 26099 25653 26111 25656
rect 26053 25647 26111 25653
rect 26970 25644 26976 25656
rect 27028 25644 27034 25696
rect 27157 25687 27215 25693
rect 27157 25653 27169 25687
rect 27203 25684 27215 25687
rect 27890 25684 27896 25696
rect 27203 25656 27896 25684
rect 27203 25653 27215 25656
rect 27157 25647 27215 25653
rect 27890 25644 27896 25656
rect 27948 25644 27954 25696
rect 36446 25644 36452 25696
rect 36504 25684 36510 25696
rect 37369 25687 37427 25693
rect 37369 25684 37381 25687
rect 36504 25656 37381 25684
rect 36504 25644 36510 25656
rect 37369 25653 37381 25656
rect 37415 25653 37427 25687
rect 37369 25647 37427 25653
rect 38105 25687 38163 25693
rect 38105 25653 38117 25687
rect 38151 25684 38163 25687
rect 38194 25684 38200 25696
rect 38151 25656 38200 25684
rect 38151 25653 38163 25656
rect 38105 25647 38163 25653
rect 38194 25644 38200 25656
rect 38252 25644 38258 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 2774 25440 2780 25492
rect 2832 25480 2838 25492
rect 9766 25480 9772 25492
rect 2832 25452 2877 25480
rect 9600 25452 9772 25480
rect 2832 25440 2838 25452
rect 6178 25304 6184 25356
rect 6236 25344 6242 25356
rect 9600 25353 9628 25452
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 11793 25483 11851 25489
rect 11793 25449 11805 25483
rect 11839 25480 11851 25483
rect 11974 25480 11980 25492
rect 11839 25452 11980 25480
rect 11839 25449 11851 25452
rect 11793 25443 11851 25449
rect 11974 25440 11980 25452
rect 12032 25440 12038 25492
rect 15010 25440 15016 25492
rect 15068 25480 15074 25492
rect 16117 25483 16175 25489
rect 16117 25480 16129 25483
rect 15068 25452 16129 25480
rect 15068 25440 15074 25452
rect 16117 25449 16129 25452
rect 16163 25449 16175 25483
rect 17402 25480 17408 25492
rect 17363 25452 17408 25480
rect 16117 25443 16175 25449
rect 6641 25347 6699 25353
rect 6641 25344 6653 25347
rect 6236 25316 6653 25344
rect 6236 25304 6242 25316
rect 6641 25313 6653 25316
rect 6687 25313 6699 25347
rect 9585 25347 9643 25353
rect 9585 25344 9597 25347
rect 6641 25307 6699 25313
rect 9048 25316 9597 25344
rect 2869 25279 2927 25285
rect 2869 25245 2881 25279
rect 2915 25276 2927 25279
rect 6546 25276 6552 25288
rect 2915 25248 6552 25276
rect 2915 25245 2927 25248
rect 2869 25239 2927 25245
rect 6546 25236 6552 25248
rect 6604 25236 6610 25288
rect 6656 25276 6684 25307
rect 9048 25276 9076 25316
rect 9585 25313 9597 25316
rect 9631 25313 9643 25347
rect 9585 25307 9643 25313
rect 11606 25304 11612 25356
rect 11664 25344 11670 25356
rect 14093 25347 14151 25353
rect 14093 25344 14105 25347
rect 11664 25316 14105 25344
rect 11664 25304 11670 25316
rect 14093 25313 14105 25316
rect 14139 25313 14151 25347
rect 14093 25307 14151 25313
rect 15102 25304 15108 25356
rect 15160 25344 15166 25356
rect 16132 25344 16160 25443
rect 17402 25440 17408 25452
rect 17460 25440 17466 25492
rect 19426 25480 19432 25492
rect 19339 25452 19432 25480
rect 19426 25440 19432 25452
rect 19484 25480 19490 25492
rect 21450 25480 21456 25492
rect 19484 25452 21456 25480
rect 19484 25440 19490 25452
rect 21450 25440 21456 25452
rect 21508 25440 21514 25492
rect 22278 25440 22284 25492
rect 22336 25480 22342 25492
rect 22373 25483 22431 25489
rect 22373 25480 22385 25483
rect 22336 25452 22385 25480
rect 22336 25440 22342 25452
rect 22373 25449 22385 25452
rect 22419 25449 22431 25483
rect 22373 25443 22431 25449
rect 22830 25440 22836 25492
rect 22888 25480 22894 25492
rect 24489 25483 24547 25489
rect 24489 25480 24501 25483
rect 22888 25452 24501 25480
rect 22888 25440 22894 25452
rect 24489 25449 24501 25452
rect 24535 25449 24547 25483
rect 25498 25480 25504 25492
rect 25459 25452 25504 25480
rect 24489 25443 24547 25449
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 25608 25452 27108 25480
rect 20257 25415 20315 25421
rect 20257 25381 20269 25415
rect 20303 25412 20315 25415
rect 20898 25412 20904 25424
rect 20303 25384 20904 25412
rect 20303 25381 20315 25384
rect 20257 25375 20315 25381
rect 20898 25372 20904 25384
rect 20956 25372 20962 25424
rect 23106 25372 23112 25424
rect 23164 25412 23170 25424
rect 25608 25412 25636 25452
rect 23164 25384 25636 25412
rect 23164 25372 23170 25384
rect 20346 25344 20352 25356
rect 15160 25316 16068 25344
rect 16132 25316 20352 25344
rect 15160 25304 15166 25316
rect 6656 25248 9076 25276
rect 9122 25236 9128 25288
rect 9180 25276 9186 25288
rect 9180 25248 9225 25276
rect 9180 25236 9186 25248
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 11882 25276 11888 25288
rect 11112 25248 11888 25276
rect 11112 25236 11118 25248
rect 11882 25236 11888 25248
rect 11940 25276 11946 25288
rect 12069 25279 12127 25285
rect 12069 25276 12081 25279
rect 11940 25248 12081 25276
rect 11940 25236 11946 25248
rect 12069 25245 12081 25248
rect 12115 25245 12127 25279
rect 12069 25239 12127 25245
rect 12161 25279 12219 25285
rect 12161 25245 12173 25279
rect 12207 25245 12219 25279
rect 12161 25239 12219 25245
rect 6908 25211 6966 25217
rect 6908 25177 6920 25211
rect 6954 25208 6966 25211
rect 7558 25208 7564 25220
rect 6954 25180 7564 25208
rect 6954 25177 6966 25180
rect 6908 25171 6966 25177
rect 7558 25168 7564 25180
rect 7616 25168 7622 25220
rect 9858 25217 9864 25220
rect 9852 25171 9864 25217
rect 9916 25208 9922 25220
rect 9916 25180 9952 25208
rect 9858 25168 9864 25171
rect 9916 25168 9922 25180
rect 8021 25143 8079 25149
rect 8021 25109 8033 25143
rect 8067 25140 8079 25143
rect 8202 25140 8208 25152
rect 8067 25112 8208 25140
rect 8067 25109 8079 25112
rect 8021 25103 8079 25109
rect 8202 25100 8208 25112
rect 8260 25100 8266 25152
rect 8478 25100 8484 25152
rect 8536 25140 8542 25152
rect 9033 25143 9091 25149
rect 9033 25140 9045 25143
rect 8536 25112 9045 25140
rect 8536 25100 8542 25112
rect 9033 25109 9045 25112
rect 9079 25109 9091 25143
rect 9033 25103 9091 25109
rect 10134 25100 10140 25152
rect 10192 25140 10198 25152
rect 10965 25143 11023 25149
rect 10965 25140 10977 25143
rect 10192 25112 10977 25140
rect 10192 25100 10198 25112
rect 10965 25109 10977 25112
rect 11011 25109 11023 25143
rect 12084 25140 12112 25239
rect 12176 25208 12204 25239
rect 12250 25236 12256 25288
rect 12308 25276 12314 25288
rect 12308 25248 12353 25276
rect 12308 25236 12314 25248
rect 12434 25236 12440 25288
rect 12492 25276 12498 25288
rect 13078 25276 13084 25288
rect 12492 25248 13084 25276
rect 12492 25236 12498 25248
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25276 13507 25279
rect 15838 25276 15844 25288
rect 13495 25248 15844 25276
rect 13495 25245 13507 25248
rect 13449 25239 13507 25245
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 16040 25276 16068 25316
rect 20346 25304 20352 25316
rect 20404 25304 20410 25356
rect 21266 25344 21272 25356
rect 21227 25316 21272 25344
rect 21266 25304 21272 25316
rect 21324 25304 21330 25356
rect 27080 25344 27108 25452
rect 27246 25440 27252 25492
rect 27304 25480 27310 25492
rect 27525 25483 27583 25489
rect 27525 25480 27537 25483
rect 27304 25452 27537 25480
rect 27304 25440 27310 25452
rect 27525 25449 27537 25452
rect 27571 25480 27583 25483
rect 28810 25480 28816 25492
rect 27571 25452 28816 25480
rect 27571 25449 27583 25452
rect 27525 25443 27583 25449
rect 28810 25440 28816 25452
rect 28868 25440 28874 25492
rect 29638 25440 29644 25492
rect 29696 25480 29702 25492
rect 29733 25483 29791 25489
rect 29733 25480 29745 25483
rect 29696 25452 29745 25480
rect 29696 25440 29702 25452
rect 29733 25449 29745 25452
rect 29779 25449 29791 25483
rect 32030 25480 32036 25492
rect 31991 25452 32036 25480
rect 29733 25443 29791 25449
rect 32030 25440 32036 25452
rect 32088 25440 32094 25492
rect 32214 25440 32220 25492
rect 32272 25480 32278 25492
rect 32769 25483 32827 25489
rect 32769 25480 32781 25483
rect 32272 25452 32781 25480
rect 32272 25440 32278 25452
rect 32769 25449 32781 25452
rect 32815 25449 32827 25483
rect 32769 25443 32827 25449
rect 29914 25344 29920 25356
rect 25976 25316 26924 25344
rect 27080 25316 28396 25344
rect 17313 25279 17371 25285
rect 16040 25248 17080 25276
rect 17052 25220 17080 25248
rect 17313 25245 17325 25279
rect 17359 25245 17371 25279
rect 17313 25239 17371 25245
rect 12342 25208 12348 25220
rect 12176 25180 12348 25208
rect 12342 25168 12348 25180
rect 12400 25168 12406 25220
rect 14360 25211 14418 25217
rect 14360 25177 14372 25211
rect 14406 25208 14418 25211
rect 14734 25208 14740 25220
rect 14406 25180 14740 25208
rect 14406 25177 14418 25180
rect 14360 25171 14418 25177
rect 14734 25168 14740 25180
rect 14792 25168 14798 25220
rect 16206 25168 16212 25220
rect 16264 25208 16270 25220
rect 16301 25211 16359 25217
rect 16301 25208 16313 25211
rect 16264 25180 16313 25208
rect 16264 25168 16270 25180
rect 16301 25177 16313 25180
rect 16347 25177 16359 25211
rect 16301 25171 16359 25177
rect 17034 25168 17040 25220
rect 17092 25208 17098 25220
rect 17328 25208 17356 25239
rect 17954 25236 17960 25288
rect 18012 25276 18018 25288
rect 18049 25279 18107 25285
rect 18049 25276 18061 25279
rect 18012 25248 18061 25276
rect 18012 25236 18018 25248
rect 18049 25245 18061 25248
rect 18095 25245 18107 25279
rect 18049 25239 18107 25245
rect 18414 25236 18420 25288
rect 18472 25276 18478 25288
rect 19242 25276 19248 25288
rect 18472 25248 19248 25276
rect 18472 25236 18478 25248
rect 19242 25236 19248 25248
rect 19300 25236 19306 25288
rect 20622 25276 20628 25288
rect 19352 25248 20628 25276
rect 19352 25208 19380 25248
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 20901 25279 20959 25285
rect 20901 25276 20913 25279
rect 20772 25248 20913 25276
rect 20772 25236 20778 25248
rect 20901 25245 20913 25248
rect 20947 25245 20959 25279
rect 22554 25276 22560 25288
rect 22467 25248 22560 25276
rect 20901 25239 20959 25245
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 22738 25276 22744 25288
rect 22699 25248 22744 25276
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 22922 25236 22928 25288
rect 22980 25276 22986 25288
rect 23293 25279 23351 25285
rect 23293 25276 23305 25279
rect 22980 25248 23305 25276
rect 22980 25236 22986 25248
rect 23293 25245 23305 25248
rect 23339 25245 23351 25279
rect 23293 25239 23351 25245
rect 23477 25279 23535 25285
rect 23477 25245 23489 25279
rect 23523 25276 23535 25279
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 23523 25248 24685 25276
rect 23523 25245 23535 25248
rect 23477 25239 23535 25245
rect 24673 25245 24685 25248
rect 24719 25276 24731 25279
rect 24762 25276 24768 25288
rect 24719 25248 24768 25276
rect 24719 25245 24731 25248
rect 24673 25239 24731 25245
rect 24762 25236 24768 25248
rect 24820 25236 24826 25288
rect 25590 25236 25596 25288
rect 25648 25276 25654 25288
rect 25976 25285 26004 25316
rect 26896 25285 26924 25316
rect 25685 25279 25743 25285
rect 25685 25276 25697 25279
rect 25648 25248 25697 25276
rect 25648 25236 25654 25248
rect 25685 25245 25697 25248
rect 25731 25245 25743 25279
rect 25685 25239 25743 25245
rect 25961 25279 26019 25285
rect 25961 25245 25973 25279
rect 26007 25245 26019 25279
rect 25961 25239 26019 25245
rect 26605 25279 26663 25285
rect 26605 25245 26617 25279
rect 26651 25245 26663 25279
rect 26605 25239 26663 25245
rect 26881 25279 26939 25285
rect 26881 25245 26893 25279
rect 26927 25276 26939 25279
rect 27062 25276 27068 25288
rect 26927 25248 27068 25276
rect 26927 25245 26939 25248
rect 26881 25239 26939 25245
rect 20070 25208 20076 25220
rect 17092 25180 19380 25208
rect 20031 25180 20076 25208
rect 17092 25168 17098 25180
rect 20070 25168 20076 25180
rect 20128 25168 20134 25220
rect 22572 25208 22600 25236
rect 22830 25208 22836 25220
rect 22572 25180 22836 25208
rect 22830 25168 22836 25180
rect 22888 25168 22894 25220
rect 25866 25208 25872 25220
rect 25779 25180 25872 25208
rect 25866 25168 25872 25180
rect 25924 25208 25930 25220
rect 26620 25208 26648 25239
rect 27062 25236 27068 25248
rect 27120 25276 27126 25288
rect 27120 25248 27568 25276
rect 27120 25236 27126 25248
rect 27540 25217 27568 25248
rect 27614 25236 27620 25288
rect 27672 25276 27678 25288
rect 28261 25279 28319 25285
rect 28261 25276 28273 25279
rect 27672 25248 28273 25276
rect 27672 25236 27678 25248
rect 28261 25245 28273 25248
rect 28307 25245 28319 25279
rect 28261 25239 28319 25245
rect 27509 25211 27568 25217
rect 25924 25180 27476 25208
rect 25924 25168 25930 25180
rect 13357 25143 13415 25149
rect 13357 25140 13369 25143
rect 12084 25112 13369 25140
rect 10965 25103 11023 25109
rect 13357 25109 13369 25112
rect 13403 25109 13415 25143
rect 15470 25140 15476 25152
rect 15431 25112 15476 25140
rect 13357 25103 13415 25109
rect 15470 25100 15476 25112
rect 15528 25100 15534 25152
rect 15746 25100 15752 25152
rect 15804 25140 15810 25152
rect 15933 25143 15991 25149
rect 15933 25140 15945 25143
rect 15804 25112 15945 25140
rect 15804 25100 15810 25112
rect 15933 25109 15945 25112
rect 15979 25109 15991 25143
rect 15933 25103 15991 25109
rect 16101 25143 16159 25149
rect 16101 25109 16113 25143
rect 16147 25140 16159 25143
rect 16574 25140 16580 25152
rect 16147 25112 16580 25140
rect 16147 25109 16159 25112
rect 16101 25103 16159 25109
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 18233 25143 18291 25149
rect 18233 25109 18245 25143
rect 18279 25140 18291 25143
rect 19150 25140 19156 25152
rect 18279 25112 19156 25140
rect 18279 25109 18291 25112
rect 18233 25103 18291 25109
rect 19150 25100 19156 25112
rect 19208 25100 19214 25152
rect 26326 25100 26332 25152
rect 26384 25140 26390 25152
rect 26421 25143 26479 25149
rect 26421 25140 26433 25143
rect 26384 25112 26433 25140
rect 26384 25100 26390 25112
rect 26421 25109 26433 25112
rect 26467 25109 26479 25143
rect 26421 25103 26479 25109
rect 26789 25143 26847 25149
rect 26789 25109 26801 25143
rect 26835 25140 26847 25143
rect 26878 25140 26884 25152
rect 26835 25112 26884 25140
rect 26835 25109 26847 25112
rect 26789 25103 26847 25109
rect 26878 25100 26884 25112
rect 26936 25100 26942 25152
rect 27338 25140 27344 25152
rect 27299 25112 27344 25140
rect 27338 25100 27344 25112
rect 27396 25100 27402 25152
rect 27448 25140 27476 25180
rect 27509 25177 27521 25211
rect 27555 25180 27568 25211
rect 27709 25211 27767 25217
rect 27709 25208 27721 25211
rect 27632 25180 27721 25208
rect 27555 25177 27567 25180
rect 27509 25171 27567 25177
rect 27632 25140 27660 25180
rect 27709 25177 27721 25180
rect 27755 25208 27767 25211
rect 27890 25208 27896 25220
rect 27755 25180 27896 25208
rect 27755 25177 27767 25180
rect 27709 25171 27767 25177
rect 27890 25168 27896 25180
rect 27948 25168 27954 25220
rect 28368 25208 28396 25316
rect 29656 25316 29920 25344
rect 29656 25285 29684 25316
rect 29914 25304 29920 25316
rect 29972 25304 29978 25356
rect 30558 25344 30564 25356
rect 30519 25316 30564 25344
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 32784 25344 32812 25443
rect 35342 25440 35348 25492
rect 35400 25480 35406 25492
rect 35437 25483 35495 25489
rect 35437 25480 35449 25483
rect 35400 25452 35449 25480
rect 35400 25440 35406 25452
rect 35437 25449 35449 25452
rect 35483 25449 35495 25483
rect 35437 25443 35495 25449
rect 33413 25415 33471 25421
rect 33413 25381 33425 25415
rect 33459 25412 33471 25415
rect 34701 25415 34759 25421
rect 34701 25412 34713 25415
rect 33459 25384 34713 25412
rect 33459 25381 33471 25384
rect 33413 25375 33471 25381
rect 34701 25381 34713 25384
rect 34747 25381 34759 25415
rect 34701 25375 34759 25381
rect 35710 25344 35716 25356
rect 32784 25316 34744 25344
rect 29641 25279 29699 25285
rect 29641 25245 29653 25279
rect 29687 25245 29699 25279
rect 29641 25239 29699 25245
rect 29825 25279 29883 25285
rect 29825 25245 29837 25279
rect 29871 25276 29883 25279
rect 30006 25276 30012 25288
rect 29871 25248 30012 25276
rect 29871 25245 29883 25248
rect 29825 25239 29883 25245
rect 30006 25236 30012 25248
rect 30064 25236 30070 25288
rect 30282 25276 30288 25288
rect 30243 25248 30288 25276
rect 30282 25236 30288 25248
rect 30340 25236 30346 25288
rect 32582 25236 32588 25288
rect 32640 25276 32646 25288
rect 32861 25279 32919 25285
rect 32861 25276 32873 25279
rect 32640 25248 32873 25276
rect 32640 25236 32646 25248
rect 32861 25245 32873 25248
rect 32907 25245 32919 25279
rect 32861 25239 32919 25245
rect 33321 25279 33379 25285
rect 33321 25245 33333 25279
rect 33367 25245 33379 25279
rect 33594 25276 33600 25288
rect 33555 25248 33600 25276
rect 33321 25239 33379 25245
rect 30834 25208 30840 25220
rect 28368 25180 30840 25208
rect 30834 25168 30840 25180
rect 30892 25168 30898 25220
rect 32490 25208 32496 25220
rect 31786 25180 32496 25208
rect 32490 25168 32496 25180
rect 32548 25168 32554 25220
rect 33336 25208 33364 25239
rect 33594 25236 33600 25248
rect 33652 25236 33658 25288
rect 34716 25285 34744 25316
rect 34900 25316 35716 25344
rect 34900 25285 34928 25316
rect 35710 25304 35716 25316
rect 35768 25304 35774 25356
rect 36262 25344 36268 25356
rect 36223 25316 36268 25344
rect 36262 25304 36268 25316
rect 36320 25304 36326 25356
rect 36446 25344 36452 25356
rect 36407 25316 36452 25344
rect 36446 25304 36452 25316
rect 36504 25304 36510 25356
rect 38102 25344 38108 25356
rect 38063 25316 38108 25344
rect 38102 25304 38108 25316
rect 38160 25304 38166 25356
rect 34701 25279 34759 25285
rect 34701 25245 34713 25279
rect 34747 25245 34759 25279
rect 34701 25239 34759 25245
rect 34885 25279 34943 25285
rect 34885 25245 34897 25279
rect 34931 25245 34943 25279
rect 35342 25276 35348 25288
rect 35303 25248 35348 25276
rect 34885 25239 34943 25245
rect 35342 25236 35348 25248
rect 35400 25236 35406 25288
rect 34054 25208 34060 25220
rect 33336 25180 34060 25208
rect 34054 25168 34060 25180
rect 34112 25168 34118 25220
rect 27448 25112 27660 25140
rect 27798 25100 27804 25152
rect 27856 25140 27862 25152
rect 28353 25143 28411 25149
rect 28353 25140 28365 25143
rect 27856 25112 28365 25140
rect 27856 25100 27862 25112
rect 28353 25109 28365 25112
rect 28399 25109 28411 25143
rect 28353 25103 28411 25109
rect 28718 25100 28724 25152
rect 28776 25140 28782 25152
rect 31202 25140 31208 25152
rect 28776 25112 31208 25140
rect 28776 25100 28782 25112
rect 31202 25100 31208 25112
rect 31260 25100 31266 25152
rect 33781 25143 33839 25149
rect 33781 25109 33793 25143
rect 33827 25140 33839 25143
rect 34606 25140 34612 25152
rect 33827 25112 34612 25140
rect 33827 25109 33839 25112
rect 33781 25103 33839 25109
rect 34606 25100 34612 25112
rect 34664 25100 34670 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 8665 24939 8723 24945
rect 8665 24905 8677 24939
rect 8711 24936 8723 24939
rect 9122 24936 9128 24948
rect 8711 24908 9128 24936
rect 8711 24905 8723 24908
rect 8665 24899 8723 24905
rect 9122 24896 9128 24908
rect 9180 24896 9186 24948
rect 11790 24896 11796 24948
rect 11848 24936 11854 24948
rect 12069 24939 12127 24945
rect 12069 24936 12081 24939
rect 11848 24908 12081 24936
rect 11848 24896 11854 24908
rect 12069 24905 12081 24908
rect 12115 24905 12127 24939
rect 14734 24936 14740 24948
rect 14695 24908 14740 24936
rect 12069 24899 12127 24905
rect 14734 24896 14740 24908
rect 14792 24896 14798 24948
rect 15105 24939 15163 24945
rect 15105 24905 15117 24939
rect 15151 24936 15163 24939
rect 15470 24936 15476 24948
rect 15151 24908 15476 24936
rect 15151 24905 15163 24908
rect 15105 24899 15163 24905
rect 15470 24896 15476 24908
rect 15528 24896 15534 24948
rect 21266 24896 21272 24948
rect 21324 24936 21330 24948
rect 25869 24939 25927 24945
rect 21324 24908 25820 24936
rect 21324 24896 21330 24908
rect 8294 24868 8300 24880
rect 8255 24840 8300 24868
rect 8294 24828 8300 24840
rect 8352 24828 8358 24880
rect 8497 24871 8555 24877
rect 8497 24868 8509 24871
rect 8496 24837 8509 24868
rect 8543 24837 8555 24871
rect 9140 24868 9168 24896
rect 12434 24868 12440 24880
rect 9140 24840 9904 24868
rect 8496 24831 8555 24837
rect 6825 24803 6883 24809
rect 6825 24769 6837 24803
rect 6871 24769 6883 24803
rect 7006 24800 7012 24812
rect 6967 24772 7012 24800
rect 6825 24763 6883 24769
rect 6840 24732 6868 24763
rect 7006 24760 7012 24772
rect 7064 24800 7070 24812
rect 7653 24803 7711 24809
rect 7653 24800 7665 24803
rect 7064 24772 7665 24800
rect 7064 24760 7070 24772
rect 7653 24769 7665 24772
rect 7699 24769 7711 24803
rect 7653 24763 7711 24769
rect 7837 24803 7895 24809
rect 7837 24769 7849 24803
rect 7883 24800 7895 24803
rect 8496 24800 8524 24831
rect 9122 24800 9128 24812
rect 7883 24772 9128 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 9122 24760 9128 24772
rect 9180 24760 9186 24812
rect 9876 24809 9904 24840
rect 11992 24840 12440 24868
rect 9769 24803 9827 24809
rect 9769 24769 9781 24803
rect 9815 24769 9827 24803
rect 9769 24763 9827 24769
rect 9861 24803 9919 24809
rect 9861 24769 9873 24803
rect 9907 24769 9919 24803
rect 9861 24763 9919 24769
rect 9953 24803 10011 24809
rect 9953 24769 9965 24803
rect 9999 24769 10011 24803
rect 10134 24800 10140 24812
rect 10095 24772 10140 24800
rect 9953 24763 10011 24769
rect 7098 24732 7104 24744
rect 6840 24704 7104 24732
rect 7098 24692 7104 24704
rect 7156 24732 7162 24744
rect 7469 24735 7527 24741
rect 7469 24732 7481 24735
rect 7156 24704 7481 24732
rect 7156 24692 7162 24704
rect 7469 24701 7481 24704
rect 7515 24701 7527 24735
rect 7469 24695 7527 24701
rect 9214 24624 9220 24676
rect 9272 24664 9278 24676
rect 9784 24664 9812 24763
rect 9968 24732 9996 24763
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 11992 24800 12020 24840
rect 12434 24828 12440 24840
rect 12492 24828 12498 24880
rect 16574 24868 16580 24880
rect 14752 24840 16580 24868
rect 11931 24772 12020 24800
rect 12161 24803 12219 24809
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12342 24800 12348 24812
rect 12207 24772 12348 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12342 24760 12348 24772
rect 12400 24800 12406 24812
rect 12805 24803 12863 24809
rect 12805 24800 12817 24803
rect 12400 24772 12817 24800
rect 12400 24760 12406 24772
rect 12805 24769 12817 24772
rect 12851 24769 12863 24803
rect 12805 24763 12863 24769
rect 13449 24803 13507 24809
rect 13449 24769 13461 24803
rect 13495 24769 13507 24803
rect 13630 24800 13636 24812
rect 13591 24772 13636 24800
rect 13449 24763 13507 24769
rect 12250 24732 12256 24744
rect 9968 24704 12256 24732
rect 12250 24692 12256 24704
rect 12308 24732 12314 24744
rect 13464 24732 13492 24763
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 13722 24760 13728 24812
rect 13780 24800 13786 24812
rect 14277 24803 14335 24809
rect 14277 24800 14289 24803
rect 13780 24772 14289 24800
rect 13780 24760 13786 24772
rect 14277 24769 14289 24772
rect 14323 24800 14335 24803
rect 14752 24800 14780 24840
rect 16574 24828 16580 24840
rect 16632 24828 16638 24880
rect 19150 24868 19156 24880
rect 19111 24840 19156 24868
rect 19150 24828 19156 24840
rect 19208 24828 19214 24880
rect 20349 24871 20407 24877
rect 20349 24837 20361 24871
rect 20395 24868 20407 24871
rect 20714 24868 20720 24880
rect 20395 24840 20720 24868
rect 20395 24837 20407 24840
rect 20349 24831 20407 24837
rect 20714 24828 20720 24840
rect 20772 24868 20778 24880
rect 20772 24840 21864 24868
rect 20772 24828 20778 24840
rect 21836 24812 21864 24840
rect 24026 24828 24032 24880
rect 24084 24828 24090 24880
rect 25792 24868 25820 24908
rect 25869 24905 25881 24939
rect 25915 24936 25927 24939
rect 27338 24936 27344 24948
rect 25915 24908 27344 24936
rect 25915 24905 25927 24908
rect 25869 24899 25927 24905
rect 27338 24896 27344 24908
rect 27396 24896 27402 24948
rect 28718 24936 28724 24948
rect 28368 24908 28724 24936
rect 28368 24868 28396 24908
rect 28718 24896 28724 24908
rect 28776 24896 28782 24948
rect 29457 24939 29515 24945
rect 29457 24905 29469 24939
rect 29503 24936 29515 24939
rect 30190 24936 30196 24948
rect 29503 24908 30196 24936
rect 29503 24905 29515 24908
rect 29457 24899 29515 24905
rect 30190 24896 30196 24908
rect 30248 24896 30254 24948
rect 30742 24896 30748 24948
rect 30800 24936 30806 24948
rect 31110 24936 31116 24948
rect 30800 24908 31116 24936
rect 30800 24896 30806 24908
rect 31110 24896 31116 24908
rect 31168 24896 31174 24948
rect 25792 24840 28396 24868
rect 28442 24828 28448 24880
rect 28500 24828 28506 24880
rect 30650 24868 30656 24880
rect 30300 24840 30656 24868
rect 14918 24800 14924 24812
rect 14323 24772 14780 24800
rect 14879 24772 14924 24800
rect 14323 24769 14335 24772
rect 14277 24763 14335 24769
rect 14918 24760 14924 24772
rect 14976 24760 14982 24812
rect 15197 24803 15255 24809
rect 15197 24769 15209 24803
rect 15243 24800 15255 24803
rect 15933 24803 15991 24809
rect 15933 24800 15945 24803
rect 15243 24772 15945 24800
rect 15243 24769 15255 24772
rect 15197 24763 15255 24769
rect 15933 24769 15945 24772
rect 15979 24769 15991 24803
rect 17034 24800 17040 24812
rect 16995 24772 17040 24800
rect 15933 24763 15991 24769
rect 12308 24704 13492 24732
rect 12308 24692 12314 24704
rect 11054 24664 11060 24676
rect 9272 24636 11060 24664
rect 9272 24624 9278 24636
rect 11054 24624 11060 24636
rect 11112 24624 11118 24676
rect 11790 24624 11796 24676
rect 11848 24664 11854 24676
rect 12713 24667 12771 24673
rect 12713 24664 12725 24667
rect 11848 24636 12725 24664
rect 11848 24624 11854 24636
rect 12713 24633 12725 24636
rect 12759 24633 12771 24667
rect 13464 24664 13492 24704
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24732 13599 24735
rect 15212 24732 15240 24763
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24800 17187 24803
rect 21177 24803 21235 24809
rect 17175 24772 18078 24800
rect 17175 24769 17187 24772
rect 17129 24763 17187 24769
rect 21177 24769 21189 24803
rect 21223 24800 21235 24803
rect 21266 24800 21272 24812
rect 21223 24772 21272 24800
rect 21223 24769 21235 24772
rect 21177 24763 21235 24769
rect 21266 24760 21272 24772
rect 21324 24800 21330 24812
rect 21634 24800 21640 24812
rect 21324 24772 21640 24800
rect 21324 24760 21330 24772
rect 21634 24760 21640 24772
rect 21692 24760 21698 24812
rect 21818 24800 21824 24812
rect 21731 24772 21824 24800
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 25961 24803 26019 24809
rect 25961 24769 25973 24803
rect 26007 24769 26019 24803
rect 27154 24800 27160 24812
rect 27115 24772 27160 24800
rect 25961 24763 26019 24769
rect 13587 24704 15240 24732
rect 13587 24701 13599 24704
rect 13541 24695 13599 24701
rect 15562 24692 15568 24744
rect 15620 24732 15626 24744
rect 15657 24735 15715 24741
rect 15657 24732 15669 24735
rect 15620 24704 15669 24732
rect 15620 24692 15626 24704
rect 15657 24701 15669 24704
rect 15703 24701 15715 24735
rect 15657 24695 15715 24701
rect 15746 24692 15752 24744
rect 15804 24732 15810 24744
rect 17681 24735 17739 24741
rect 15804 24704 15849 24732
rect 15804 24692 15810 24704
rect 17681 24701 17693 24735
rect 17727 24732 17739 24735
rect 18506 24732 18512 24744
rect 17727 24704 18512 24732
rect 17727 24701 17739 24704
rect 17681 24695 17739 24701
rect 18506 24692 18512 24704
rect 18564 24692 18570 24744
rect 19429 24735 19487 24741
rect 19429 24732 19441 24735
rect 19352 24704 19441 24732
rect 14458 24664 14464 24676
rect 13464 24636 14464 24664
rect 12713 24627 12771 24633
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 6914 24596 6920 24608
rect 6875 24568 6920 24596
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 8202 24556 8208 24608
rect 8260 24596 8266 24608
rect 8481 24599 8539 24605
rect 8481 24596 8493 24599
rect 8260 24568 8493 24596
rect 8260 24556 8266 24568
rect 8481 24565 8493 24568
rect 8527 24565 8539 24599
rect 8481 24559 8539 24565
rect 9493 24599 9551 24605
rect 9493 24565 9505 24599
rect 9539 24596 9551 24599
rect 9766 24596 9772 24608
rect 9539 24568 9772 24596
rect 9539 24565 9551 24568
rect 9493 24559 9551 24565
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 11885 24599 11943 24605
rect 11885 24565 11897 24599
rect 11931 24596 11943 24599
rect 12158 24596 12164 24608
rect 11931 24568 12164 24596
rect 11931 24565 11943 24568
rect 11885 24559 11943 24565
rect 12158 24556 12164 24568
rect 12216 24556 12222 24608
rect 14182 24596 14188 24608
rect 14143 24568 14188 24596
rect 14182 24556 14188 24568
rect 14240 24556 14246 24608
rect 16114 24596 16120 24608
rect 16075 24568 16120 24596
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 19352 24596 19380 24704
rect 19429 24701 19441 24704
rect 19475 24701 19487 24735
rect 19429 24695 19487 24701
rect 22094 24692 22100 24744
rect 22152 24732 22158 24744
rect 22152 24704 22197 24732
rect 22152 24692 22158 24704
rect 23198 24692 23204 24744
rect 23256 24732 23262 24744
rect 23293 24735 23351 24741
rect 23293 24732 23305 24735
rect 23256 24704 23305 24732
rect 23256 24692 23262 24704
rect 23293 24701 23305 24704
rect 23339 24701 23351 24735
rect 23566 24732 23572 24744
rect 23527 24704 23572 24732
rect 23293 24695 23351 24701
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24701 25099 24735
rect 25041 24695 25099 24701
rect 25056 24664 25084 24695
rect 25406 24692 25412 24744
rect 25464 24732 25470 24744
rect 25976 24732 26004 24763
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 29730 24760 29736 24812
rect 29788 24800 29794 24812
rect 30009 24803 30067 24809
rect 30009 24800 30021 24803
rect 29788 24772 30021 24800
rect 29788 24760 29794 24772
rect 30009 24769 30021 24772
rect 30055 24769 30067 24803
rect 30009 24763 30067 24769
rect 30193 24803 30251 24809
rect 30193 24769 30205 24803
rect 30239 24800 30251 24803
rect 30300 24800 30328 24840
rect 30650 24828 30656 24840
rect 30708 24828 30714 24880
rect 31570 24868 31576 24880
rect 30852 24840 31576 24868
rect 30239 24772 30328 24800
rect 30239 24769 30251 24772
rect 30193 24763 30251 24769
rect 30374 24760 30380 24812
rect 30432 24800 30438 24812
rect 30852 24809 30880 24840
rect 31570 24828 31576 24840
rect 31628 24828 31634 24880
rect 30837 24803 30895 24809
rect 30432 24772 30477 24800
rect 30432 24760 30438 24772
rect 30837 24769 30849 24803
rect 30883 24769 30895 24803
rect 30837 24763 30895 24769
rect 30926 24760 30932 24812
rect 30984 24800 30990 24812
rect 31110 24800 31116 24812
rect 30984 24772 31029 24800
rect 31071 24772 31116 24800
rect 30984 24760 30990 24772
rect 31110 24760 31116 24772
rect 31168 24760 31174 24812
rect 33502 24760 33508 24812
rect 33560 24760 33566 24812
rect 34330 24800 34336 24812
rect 33612 24772 33992 24800
rect 34291 24772 34336 24800
rect 25464 24704 26004 24732
rect 25464 24692 25470 24704
rect 26142 24692 26148 24744
rect 26200 24732 26206 24744
rect 27706 24732 27712 24744
rect 26200 24704 26245 24732
rect 26344 24704 27712 24732
rect 26200 24692 26206 24704
rect 25958 24664 25964 24676
rect 25056 24636 25964 24664
rect 25958 24624 25964 24636
rect 26016 24624 26022 24676
rect 26344 24664 26372 24704
rect 27706 24692 27712 24704
rect 27764 24692 27770 24744
rect 27985 24735 28043 24741
rect 27985 24701 27997 24735
rect 28031 24732 28043 24735
rect 28350 24732 28356 24744
rect 28031 24704 28356 24732
rect 28031 24701 28043 24704
rect 27985 24695 28043 24701
rect 28350 24692 28356 24704
rect 28408 24692 28414 24744
rect 30282 24692 30288 24744
rect 30340 24732 30346 24744
rect 32125 24735 32183 24741
rect 32125 24732 32137 24735
rect 30340 24704 32137 24732
rect 30340 24692 30346 24704
rect 32125 24701 32137 24704
rect 32171 24701 32183 24735
rect 32398 24732 32404 24744
rect 32359 24704 32404 24732
rect 32125 24695 32183 24701
rect 26160 24636 26372 24664
rect 26160 24608 26188 24636
rect 26694 24624 26700 24676
rect 26752 24664 26758 24676
rect 26752 24636 27108 24664
rect 26752 24624 26758 24636
rect 17920 24568 19380 24596
rect 17920 24556 17926 24568
rect 25130 24556 25136 24608
rect 25188 24596 25194 24608
rect 25501 24599 25559 24605
rect 25501 24596 25513 24599
rect 25188 24568 25513 24596
rect 25188 24556 25194 24568
rect 25501 24565 25513 24568
rect 25547 24565 25559 24599
rect 25501 24559 25559 24565
rect 26142 24556 26148 24608
rect 26200 24556 26206 24608
rect 26418 24556 26424 24608
rect 26476 24596 26482 24608
rect 26973 24599 27031 24605
rect 26973 24596 26985 24599
rect 26476 24568 26985 24596
rect 26476 24556 26482 24568
rect 26973 24565 26985 24568
rect 27019 24565 27031 24599
rect 27080 24596 27108 24636
rect 30466 24624 30472 24676
rect 30524 24664 30530 24676
rect 30837 24667 30895 24673
rect 30837 24664 30849 24667
rect 30524 24636 30849 24664
rect 30524 24624 30530 24636
rect 30837 24633 30849 24636
rect 30883 24633 30895 24667
rect 30837 24627 30895 24633
rect 31386 24596 31392 24608
rect 27080 24568 31392 24596
rect 26973 24559 27031 24565
rect 31386 24556 31392 24568
rect 31444 24556 31450 24608
rect 32030 24556 32036 24608
rect 32088 24596 32094 24608
rect 32140 24596 32168 24695
rect 32398 24692 32404 24704
rect 32456 24692 32462 24744
rect 32950 24692 32956 24744
rect 33008 24732 33014 24744
rect 33612 24732 33640 24772
rect 33008 24704 33640 24732
rect 33008 24692 33014 24704
rect 33778 24692 33784 24744
rect 33836 24732 33842 24744
rect 33873 24735 33931 24741
rect 33873 24732 33885 24735
rect 33836 24704 33885 24732
rect 33836 24692 33842 24704
rect 33873 24701 33885 24704
rect 33919 24701 33931 24735
rect 33964 24732 33992 24772
rect 34330 24760 34336 24772
rect 34388 24760 34394 24812
rect 35710 24760 35716 24812
rect 35768 24760 35774 24812
rect 34606 24732 34612 24744
rect 33964 24704 34468 24732
rect 34567 24704 34612 24732
rect 33873 24695 33931 24701
rect 34330 24664 34336 24676
rect 33428 24636 34336 24664
rect 33428 24596 33456 24636
rect 34330 24624 34336 24636
rect 34388 24624 34394 24676
rect 32088 24568 33456 24596
rect 34440 24596 34468 24704
rect 34606 24692 34612 24704
rect 34664 24692 34670 24744
rect 35802 24692 35808 24744
rect 35860 24732 35866 24744
rect 36081 24735 36139 24741
rect 36081 24732 36093 24735
rect 35860 24704 36093 24732
rect 35860 24692 35866 24704
rect 36081 24701 36093 24704
rect 36127 24701 36139 24735
rect 36081 24695 36139 24701
rect 37274 24664 37280 24676
rect 35636 24636 37280 24664
rect 35636 24596 35664 24636
rect 37274 24624 37280 24636
rect 37332 24624 37338 24676
rect 34440 24568 35664 24596
rect 32088 24556 32094 24568
rect 36262 24556 36268 24608
rect 36320 24596 36326 24608
rect 36541 24599 36599 24605
rect 36541 24596 36553 24599
rect 36320 24568 36553 24596
rect 36320 24556 36326 24568
rect 36541 24565 36553 24568
rect 36587 24565 36599 24599
rect 37826 24596 37832 24608
rect 37787 24568 37832 24596
rect 36541 24559 36599 24565
rect 37826 24556 37832 24568
rect 37884 24556 37890 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 7558 24392 7564 24404
rect 7519 24364 7564 24392
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 9122 24392 9128 24404
rect 9083 24364 9128 24392
rect 9122 24352 9128 24364
rect 9180 24352 9186 24404
rect 9858 24392 9864 24404
rect 9819 24364 9864 24392
rect 9858 24352 9864 24364
rect 9916 24352 9922 24404
rect 13081 24395 13139 24401
rect 13081 24361 13093 24395
rect 13127 24392 13139 24395
rect 14090 24392 14096 24404
rect 13127 24364 14096 24392
rect 13127 24361 13139 24364
rect 13081 24355 13139 24361
rect 14090 24352 14096 24364
rect 14148 24352 14154 24404
rect 14918 24392 14924 24404
rect 14879 24364 14924 24392
rect 14918 24352 14924 24364
rect 14976 24352 14982 24404
rect 15105 24395 15163 24401
rect 15105 24361 15117 24395
rect 15151 24392 15163 24395
rect 15562 24392 15568 24404
rect 15151 24364 15568 24392
rect 15151 24361 15163 24364
rect 15105 24355 15163 24361
rect 15562 24352 15568 24364
rect 15620 24352 15626 24404
rect 18322 24352 18328 24404
rect 18380 24392 18386 24404
rect 18601 24395 18659 24401
rect 18601 24392 18613 24395
rect 18380 24364 18613 24392
rect 18380 24352 18386 24364
rect 18601 24361 18613 24364
rect 18647 24392 18659 24395
rect 18647 24364 23244 24392
rect 18647 24361 18659 24364
rect 18601 24355 18659 24361
rect 8294 24284 8300 24336
rect 8352 24324 8358 24336
rect 13265 24327 13323 24333
rect 8352 24296 8984 24324
rect 8352 24284 8358 24296
rect 8478 24256 8484 24268
rect 7852 24228 8484 24256
rect 7006 24188 7012 24200
rect 6967 24160 7012 24188
rect 7006 24148 7012 24160
rect 7064 24148 7070 24200
rect 7650 24148 7656 24200
rect 7708 24188 7714 24200
rect 7852 24197 7880 24228
rect 8478 24216 8484 24228
rect 8536 24216 8542 24268
rect 8956 24265 8984 24296
rect 13265 24293 13277 24327
rect 13311 24324 13323 24327
rect 13722 24324 13728 24336
rect 13311 24296 13728 24324
rect 13311 24293 13323 24296
rect 13265 24287 13323 24293
rect 13722 24284 13728 24296
rect 13780 24284 13786 24336
rect 14185 24327 14243 24333
rect 14185 24293 14197 24327
rect 14231 24324 14243 24327
rect 14274 24324 14280 24336
rect 14231 24296 14280 24324
rect 14231 24293 14243 24296
rect 14185 24287 14243 24293
rect 14274 24284 14280 24296
rect 14332 24324 14338 24336
rect 16298 24324 16304 24336
rect 14332 24296 16304 24324
rect 14332 24284 14338 24296
rect 16298 24284 16304 24296
rect 16356 24284 16362 24336
rect 17865 24327 17923 24333
rect 17865 24293 17877 24327
rect 17911 24324 17923 24327
rect 20441 24327 20499 24333
rect 17911 24296 20392 24324
rect 17911 24293 17923 24296
rect 17865 24287 17923 24293
rect 8941 24259 8999 24265
rect 8941 24225 8953 24259
rect 8987 24225 8999 24259
rect 15470 24256 15476 24268
rect 15431 24228 15476 24256
rect 8941 24219 8999 24225
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 20364 24256 20392 24296
rect 20441 24293 20453 24327
rect 20487 24324 20499 24327
rect 22922 24324 22928 24336
rect 20487 24296 22928 24324
rect 20487 24293 20499 24296
rect 20441 24287 20499 24293
rect 22922 24284 22928 24296
rect 22980 24284 22986 24336
rect 21174 24256 21180 24268
rect 17972 24228 20300 24256
rect 20364 24228 21180 24256
rect 7745 24191 7803 24197
rect 7745 24188 7757 24191
rect 7708 24160 7757 24188
rect 7708 24148 7714 24160
rect 7745 24157 7757 24160
rect 7791 24157 7803 24191
rect 7745 24151 7803 24157
rect 7837 24191 7895 24197
rect 7837 24157 7849 24191
rect 7883 24157 7895 24191
rect 8202 24188 8208 24200
rect 8163 24160 8208 24188
rect 7837 24151 7895 24157
rect 8202 24148 8208 24160
rect 8260 24148 8266 24200
rect 9214 24188 9220 24200
rect 9175 24160 9220 24188
rect 9214 24148 9220 24160
rect 9272 24148 9278 24200
rect 9674 24188 9680 24200
rect 9635 24160 9680 24188
rect 9674 24148 9680 24160
rect 9732 24148 9738 24200
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 9861 24191 9919 24197
rect 9861 24188 9873 24191
rect 9824 24160 9873 24188
rect 9824 24148 9830 24160
rect 9861 24157 9873 24160
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24188 10655 24191
rect 11606 24188 11612 24200
rect 10643 24160 11612 24188
rect 10643 24157 10655 24160
rect 10597 24151 10655 24157
rect 11606 24148 11612 24160
rect 11664 24148 11670 24200
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 12308 24160 13032 24188
rect 12308 24148 12314 24160
rect 6825 24123 6883 24129
rect 6825 24089 6837 24123
rect 6871 24120 6883 24123
rect 7098 24120 7104 24132
rect 6871 24092 7104 24120
rect 6871 24089 6883 24092
rect 6825 24083 6883 24089
rect 7098 24080 7104 24092
rect 7156 24080 7162 24132
rect 7929 24123 7987 24129
rect 7929 24089 7941 24123
rect 7975 24089 7987 24123
rect 7929 24083 7987 24089
rect 8067 24123 8125 24129
rect 8067 24089 8079 24123
rect 8113 24120 8125 24123
rect 9490 24120 9496 24132
rect 8113 24092 9496 24120
rect 8113 24089 8125 24092
rect 8067 24083 8125 24089
rect 6546 24012 6552 24064
rect 6604 24052 6610 24064
rect 6641 24055 6699 24061
rect 6641 24052 6653 24055
rect 6604 24024 6653 24052
rect 6604 24012 6610 24024
rect 6641 24021 6653 24024
rect 6687 24021 6699 24055
rect 7944 24052 7972 24083
rect 9490 24080 9496 24092
rect 9548 24080 9554 24132
rect 10864 24123 10922 24129
rect 10864 24089 10876 24123
rect 10910 24120 10922 24123
rect 11514 24120 11520 24132
rect 10910 24092 11520 24120
rect 10910 24089 10922 24092
rect 10864 24083 10922 24089
rect 11514 24080 11520 24092
rect 11572 24080 11578 24132
rect 12434 24080 12440 24132
rect 12492 24120 12498 24132
rect 12897 24123 12955 24129
rect 12897 24120 12909 24123
rect 12492 24092 12909 24120
rect 12492 24080 12498 24092
rect 12897 24089 12909 24092
rect 12943 24089 12955 24123
rect 13004 24120 13032 24160
rect 16666 24148 16672 24200
rect 16724 24188 16730 24200
rect 17310 24188 17316 24200
rect 16724 24160 17316 24188
rect 16724 24148 16730 24160
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 17972 24197 18000 24228
rect 17957 24191 18015 24197
rect 17957 24157 17969 24191
rect 18003 24157 18015 24191
rect 17957 24151 18015 24157
rect 18417 24191 18475 24197
rect 18417 24157 18429 24191
rect 18463 24188 18475 24191
rect 19242 24188 19248 24200
rect 18463 24160 19248 24188
rect 18463 24157 18475 24160
rect 18417 24151 18475 24157
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 13097 24123 13155 24129
rect 13097 24120 13109 24123
rect 13004 24092 13109 24120
rect 12897 24083 12955 24089
rect 13097 24089 13109 24092
rect 13143 24089 13155 24123
rect 14366 24120 14372 24132
rect 14327 24092 14372 24120
rect 13097 24083 13155 24089
rect 14366 24080 14372 24092
rect 14424 24080 14430 24132
rect 15105 24123 15163 24129
rect 15105 24089 15117 24123
rect 15151 24120 15163 24123
rect 15746 24120 15752 24132
rect 15151 24092 15752 24120
rect 15151 24089 15163 24092
rect 15105 24083 15163 24089
rect 15746 24080 15752 24092
rect 15804 24080 15810 24132
rect 16114 24080 16120 24132
rect 16172 24120 16178 24132
rect 17046 24123 17104 24129
rect 17046 24120 17058 24123
rect 16172 24092 17058 24120
rect 16172 24080 16178 24092
rect 17046 24089 17058 24092
rect 17092 24089 17104 24123
rect 17046 24083 17104 24089
rect 19429 24123 19487 24129
rect 19429 24089 19441 24123
rect 19475 24120 19487 24123
rect 20162 24120 20168 24132
rect 19475 24092 20168 24120
rect 19475 24089 19487 24092
rect 19429 24083 19487 24089
rect 20162 24080 20168 24092
rect 20220 24080 20226 24132
rect 20272 24129 20300 24228
rect 21174 24216 21180 24228
rect 21232 24216 21238 24268
rect 21545 24259 21603 24265
rect 21545 24225 21557 24259
rect 21591 24225 21603 24259
rect 23216 24256 23244 24364
rect 23566 24352 23572 24404
rect 23624 24392 23630 24404
rect 24397 24395 24455 24401
rect 24397 24392 24409 24395
rect 23624 24364 24409 24392
rect 23624 24352 23630 24364
rect 24397 24361 24409 24364
rect 24443 24361 24455 24395
rect 24397 24355 24455 24361
rect 25685 24395 25743 24401
rect 25685 24361 25697 24395
rect 25731 24392 25743 24395
rect 27154 24392 27160 24404
rect 25731 24364 27160 24392
rect 25731 24361 25743 24364
rect 25685 24355 25743 24361
rect 27154 24352 27160 24364
rect 27212 24352 27218 24404
rect 27890 24392 27896 24404
rect 27851 24364 27896 24392
rect 27890 24352 27896 24364
rect 27948 24352 27954 24404
rect 28350 24392 28356 24404
rect 28311 24364 28356 24392
rect 28350 24352 28356 24364
rect 28408 24352 28414 24404
rect 32490 24392 32496 24404
rect 28966 24364 31754 24392
rect 32451 24364 32496 24392
rect 23753 24327 23811 24333
rect 23753 24293 23765 24327
rect 23799 24324 23811 24327
rect 24026 24324 24032 24336
rect 23799 24296 24032 24324
rect 23799 24293 23811 24296
rect 23753 24287 23811 24293
rect 24026 24284 24032 24296
rect 24084 24284 24090 24336
rect 25774 24256 25780 24268
rect 23216 24228 25780 24256
rect 21545 24219 21603 24225
rect 20257 24123 20315 24129
rect 20257 24089 20269 24123
rect 20303 24120 20315 24123
rect 20622 24120 20628 24132
rect 20303 24092 20628 24120
rect 20303 24089 20315 24092
rect 20257 24083 20315 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 8478 24052 8484 24064
rect 7944 24024 8484 24052
rect 6641 24015 6699 24021
rect 8478 24012 8484 24024
rect 8536 24012 8542 24064
rect 8570 24012 8576 24064
rect 8628 24052 8634 24064
rect 8941 24055 8999 24061
rect 8941 24052 8953 24055
rect 8628 24024 8953 24052
rect 8628 24012 8634 24024
rect 8941 24021 8953 24024
rect 8987 24021 8999 24055
rect 9508 24052 9536 24080
rect 11882 24052 11888 24064
rect 9508 24024 11888 24052
rect 8941 24015 8999 24021
rect 11882 24012 11888 24024
rect 11940 24012 11946 24064
rect 11977 24055 12035 24061
rect 11977 24021 11989 24055
rect 12023 24052 12035 24055
rect 12158 24052 12164 24064
rect 12023 24024 12164 24052
rect 12023 24021 12035 24024
rect 11977 24015 12035 24021
rect 12158 24012 12164 24024
rect 12216 24012 12222 24064
rect 15562 24012 15568 24064
rect 15620 24052 15626 24064
rect 15933 24055 15991 24061
rect 15933 24052 15945 24055
rect 15620 24024 15945 24052
rect 15620 24012 15626 24024
rect 15933 24021 15945 24024
rect 15979 24021 15991 24055
rect 15933 24015 15991 24021
rect 17770 24012 17776 24064
rect 17828 24052 17834 24064
rect 20990 24052 20996 24064
rect 17828 24024 20996 24052
rect 17828 24012 17834 24024
rect 20990 24012 20996 24024
rect 21048 24052 21054 24064
rect 21560 24052 21588 24219
rect 25774 24216 25780 24228
rect 25832 24216 25838 24268
rect 26418 24256 26424 24268
rect 26379 24228 26424 24256
rect 26418 24216 26424 24228
rect 26476 24216 26482 24268
rect 21818 24188 21824 24200
rect 21779 24160 21824 24188
rect 21818 24148 21824 24160
rect 21876 24188 21882 24200
rect 22465 24191 22523 24197
rect 22465 24188 22477 24191
rect 21876 24160 22477 24188
rect 21876 24148 21882 24160
rect 22465 24157 22477 24160
rect 22511 24157 22523 24191
rect 23658 24188 23664 24200
rect 23619 24160 23664 24188
rect 22465 24151 22523 24157
rect 23658 24148 23664 24160
rect 23716 24148 23722 24200
rect 24581 24191 24639 24197
rect 24581 24157 24593 24191
rect 24627 24188 24639 24191
rect 25130 24188 25136 24200
rect 24627 24160 25136 24188
rect 24627 24157 24639 24160
rect 24581 24151 24639 24157
rect 25130 24148 25136 24160
rect 25188 24148 25194 24200
rect 25406 24188 25412 24200
rect 25367 24160 25412 24188
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 25501 24191 25559 24197
rect 25501 24157 25513 24191
rect 25547 24157 25559 24191
rect 26142 24188 26148 24200
rect 26103 24160 26148 24188
rect 25501 24151 25559 24157
rect 23014 24080 23020 24132
rect 23072 24120 23078 24132
rect 25516 24120 25544 24151
rect 26142 24148 26148 24160
rect 26200 24148 26206 24200
rect 28534 24188 28540 24200
rect 28495 24160 28540 24188
rect 28534 24148 28540 24160
rect 28592 24148 28598 24200
rect 26326 24120 26332 24132
rect 23072 24092 23117 24120
rect 25516 24092 26332 24120
rect 23072 24080 23078 24092
rect 26326 24080 26332 24092
rect 26384 24080 26390 24132
rect 27430 24080 27436 24132
rect 27488 24080 27494 24132
rect 28966 24052 28994 24364
rect 31726 24324 31754 24364
rect 32490 24352 32496 24364
rect 32548 24352 32554 24404
rect 33137 24395 33195 24401
rect 33137 24361 33149 24395
rect 33183 24392 33195 24395
rect 33502 24392 33508 24404
rect 33183 24364 33508 24392
rect 33183 24361 33195 24364
rect 33137 24355 33195 24361
rect 33502 24352 33508 24364
rect 33560 24352 33566 24404
rect 34793 24395 34851 24401
rect 34793 24361 34805 24395
rect 34839 24392 34851 24395
rect 35710 24392 35716 24404
rect 34839 24364 35716 24392
rect 34839 24361 34851 24364
rect 34793 24355 34851 24361
rect 35710 24352 35716 24364
rect 35768 24352 35774 24404
rect 32950 24324 32956 24336
rect 31726 24296 32956 24324
rect 32950 24284 32956 24296
rect 33008 24284 33014 24336
rect 34698 24324 34704 24336
rect 33060 24296 34704 24324
rect 29546 24256 29552 24268
rect 29459 24228 29552 24256
rect 29546 24216 29552 24228
rect 29604 24256 29610 24268
rect 30282 24256 30288 24268
rect 29604 24228 30288 24256
rect 29604 24216 29610 24228
rect 30282 24216 30288 24228
rect 30340 24216 30346 24268
rect 31938 24188 31944 24200
rect 31851 24160 31944 24188
rect 31938 24148 31944 24160
rect 31996 24188 32002 24200
rect 33060 24197 33088 24296
rect 34698 24284 34704 24296
rect 34756 24284 34762 24336
rect 33502 24216 33508 24268
rect 33560 24256 33566 24268
rect 36262 24256 36268 24268
rect 33560 24228 35480 24256
rect 36223 24228 36268 24256
rect 33560 24216 33566 24228
rect 35452 24200 35480 24228
rect 36262 24216 36268 24228
rect 36320 24216 36326 24268
rect 32585 24191 32643 24197
rect 32585 24188 32597 24191
rect 31996 24160 32597 24188
rect 31996 24148 32002 24160
rect 32585 24157 32597 24160
rect 32631 24188 32643 24191
rect 33045 24191 33103 24197
rect 33045 24188 33057 24191
rect 32631 24160 33057 24188
rect 32631 24157 32643 24160
rect 32585 24151 32643 24157
rect 33045 24157 33057 24160
rect 33091 24157 33103 24191
rect 33045 24151 33103 24157
rect 34149 24191 34207 24197
rect 34149 24157 34161 24191
rect 34195 24188 34207 24191
rect 34606 24188 34612 24200
rect 34195 24160 34612 24188
rect 34195 24157 34207 24160
rect 34149 24151 34207 24157
rect 34606 24148 34612 24160
rect 34664 24148 34670 24200
rect 34698 24148 34704 24200
rect 34756 24188 34762 24200
rect 35342 24188 35348 24200
rect 34756 24160 35348 24188
rect 34756 24148 34762 24160
rect 35342 24148 35348 24160
rect 35400 24148 35406 24200
rect 35434 24148 35440 24200
rect 35492 24188 35498 24200
rect 35529 24191 35587 24197
rect 35529 24188 35541 24191
rect 35492 24160 35541 24188
rect 35492 24148 35498 24160
rect 35529 24157 35541 24160
rect 35575 24157 35587 24191
rect 35529 24151 35587 24157
rect 29822 24120 29828 24132
rect 29783 24092 29828 24120
rect 29822 24080 29828 24092
rect 29880 24080 29886 24132
rect 31849 24123 31907 24129
rect 31849 24120 31861 24123
rect 31050 24092 31861 24120
rect 31849 24089 31861 24092
rect 31895 24089 31907 24123
rect 31849 24083 31907 24089
rect 32766 24080 32772 24132
rect 32824 24120 32830 24132
rect 34422 24120 34428 24132
rect 32824 24092 34428 24120
rect 32824 24080 32830 24092
rect 34422 24080 34428 24092
rect 34480 24080 34486 24132
rect 34514 24080 34520 24132
rect 34572 24120 34578 24132
rect 36449 24123 36507 24129
rect 34572 24092 35572 24120
rect 34572 24080 34578 24092
rect 35544 24064 35572 24092
rect 36449 24089 36461 24123
rect 36495 24120 36507 24123
rect 37366 24120 37372 24132
rect 36495 24092 37372 24120
rect 36495 24089 36507 24092
rect 36449 24083 36507 24089
rect 37366 24080 37372 24092
rect 37424 24080 37430 24132
rect 38102 24120 38108 24132
rect 38063 24092 38108 24120
rect 38102 24080 38108 24092
rect 38160 24080 38166 24132
rect 21048 24024 28994 24052
rect 21048 24012 21054 24024
rect 30650 24012 30656 24064
rect 30708 24052 30714 24064
rect 31297 24055 31355 24061
rect 31297 24052 31309 24055
rect 30708 24024 31309 24052
rect 30708 24012 30714 24024
rect 31297 24021 31309 24024
rect 31343 24021 31355 24055
rect 31297 24015 31355 24021
rect 31386 24012 31392 24064
rect 31444 24052 31450 24064
rect 34882 24052 34888 24064
rect 31444 24024 34888 24052
rect 31444 24012 31450 24024
rect 34882 24012 34888 24024
rect 34940 24012 34946 24064
rect 35342 24012 35348 24064
rect 35400 24052 35406 24064
rect 35437 24055 35495 24061
rect 35437 24052 35449 24055
rect 35400 24024 35449 24052
rect 35400 24012 35406 24024
rect 35437 24021 35449 24024
rect 35483 24021 35495 24055
rect 35437 24015 35495 24021
rect 35526 24012 35532 24064
rect 35584 24012 35590 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 6914 23808 6920 23860
rect 6972 23808 6978 23860
rect 7650 23848 7656 23860
rect 7611 23820 7656 23848
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 8294 23848 8300 23860
rect 7944 23820 8300 23848
rect 6733 23783 6791 23789
rect 6733 23749 6745 23783
rect 6779 23780 6791 23783
rect 6932 23780 6960 23808
rect 6779 23752 6960 23780
rect 6779 23749 6791 23752
rect 6733 23743 6791 23749
rect 7006 23740 7012 23792
rect 7064 23780 7070 23792
rect 7742 23780 7748 23792
rect 7064 23752 7748 23780
rect 7064 23740 7070 23752
rect 7742 23740 7748 23752
rect 7800 23780 7806 23792
rect 7800 23752 7880 23780
rect 7800 23740 7806 23752
rect 6546 23712 6552 23724
rect 6507 23684 6552 23712
rect 6546 23672 6552 23684
rect 6604 23672 6610 23724
rect 6638 23672 6644 23724
rect 6696 23712 6702 23724
rect 7852 23721 7880 23752
rect 7944 23721 7972 23820
rect 8294 23808 8300 23820
rect 8352 23848 8358 23860
rect 10229 23851 10287 23857
rect 10229 23848 10241 23851
rect 8352 23820 10241 23848
rect 8352 23808 8358 23820
rect 10229 23817 10241 23820
rect 10275 23817 10287 23851
rect 11514 23848 11520 23860
rect 11475 23820 11520 23848
rect 10229 23811 10287 23817
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 11882 23808 11888 23860
rect 11940 23848 11946 23860
rect 13354 23848 13360 23860
rect 11940 23820 13360 23848
rect 11940 23808 11946 23820
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 13630 23808 13636 23860
rect 13688 23848 13694 23860
rect 15105 23851 15163 23857
rect 15105 23848 15117 23851
rect 13688 23820 15117 23848
rect 13688 23808 13694 23820
rect 15105 23817 15117 23820
rect 15151 23817 15163 23851
rect 15105 23811 15163 23817
rect 19981 23851 20039 23857
rect 19981 23817 19993 23851
rect 20027 23848 20039 23851
rect 20070 23848 20076 23860
rect 20027 23820 20076 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 20070 23808 20076 23820
rect 20128 23808 20134 23860
rect 22094 23808 22100 23860
rect 22152 23848 22158 23860
rect 23750 23848 23756 23860
rect 22152 23820 23756 23848
rect 22152 23808 22158 23820
rect 23750 23808 23756 23820
rect 23808 23808 23814 23860
rect 24118 23848 24124 23860
rect 24079 23820 24124 23848
rect 24118 23808 24124 23820
rect 24176 23808 24182 23860
rect 24489 23851 24547 23857
rect 24489 23817 24501 23851
rect 24535 23848 24547 23851
rect 24670 23848 24676 23860
rect 24535 23820 24676 23848
rect 24535 23817 24547 23820
rect 24489 23811 24547 23817
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 25409 23851 25467 23857
rect 25409 23817 25421 23851
rect 25455 23848 25467 23851
rect 27246 23848 27252 23860
rect 25455 23820 27252 23848
rect 25455 23817 25467 23820
rect 25409 23811 25467 23817
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 27341 23851 27399 23857
rect 27341 23817 27353 23851
rect 27387 23848 27399 23851
rect 27430 23848 27436 23860
rect 27387 23820 27436 23848
rect 27387 23817 27399 23820
rect 27341 23811 27399 23817
rect 27430 23808 27436 23820
rect 27488 23808 27494 23860
rect 32766 23848 32772 23860
rect 31726 23820 32772 23848
rect 8202 23780 8208 23792
rect 8115 23752 8208 23780
rect 8128 23721 8156 23752
rect 8202 23740 8208 23752
rect 8260 23780 8266 23792
rect 8260 23752 9628 23780
rect 8260 23740 8266 23752
rect 6851 23715 6909 23721
rect 6851 23712 6863 23715
rect 6696 23684 6741 23712
rect 6696 23672 6702 23684
rect 6840 23681 6863 23712
rect 6897 23681 6909 23715
rect 6840 23675 6909 23681
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23681 7895 23715
rect 7837 23675 7895 23681
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 8113 23715 8171 23721
rect 8113 23681 8125 23715
rect 8159 23681 8171 23715
rect 8846 23712 8852 23724
rect 8807 23684 8852 23712
rect 8113 23675 8171 23681
rect 6840 23644 6868 23675
rect 8846 23672 8852 23684
rect 8904 23672 8910 23724
rect 9600 23721 9628 23752
rect 11606 23740 11612 23792
rect 11664 23780 11670 23792
rect 11664 23752 12434 23780
rect 11664 23740 11670 23752
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23712 9643 23715
rect 9674 23712 9680 23724
rect 9631 23684 9680 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 9674 23672 9680 23684
rect 9732 23672 9738 23724
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23712 9827 23715
rect 10134 23712 10140 23724
rect 9815 23684 10140 23712
rect 9815 23681 9827 23684
rect 9769 23675 9827 23681
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 10410 23712 10416 23724
rect 10371 23684 10416 23712
rect 10410 23672 10416 23684
rect 10468 23672 10474 23724
rect 11701 23715 11759 23721
rect 11701 23681 11713 23715
rect 11747 23681 11759 23715
rect 11793 23715 11851 23721
rect 11793 23708 11805 23715
rect 11839 23708 11851 23715
rect 11885 23715 11943 23721
rect 11701 23675 11759 23681
rect 6748 23616 6868 23644
rect 7009 23647 7067 23653
rect 6748 23588 6776 23616
rect 7009 23613 7021 23647
rect 7055 23644 7067 23647
rect 7098 23644 7104 23656
rect 7055 23616 7104 23644
rect 7055 23613 7067 23616
rect 7009 23607 7067 23613
rect 7098 23604 7104 23616
rect 7156 23644 7162 23656
rect 8021 23647 8079 23653
rect 8021 23644 8033 23647
rect 7156 23616 8033 23644
rect 7156 23604 7162 23616
rect 8021 23613 8033 23616
rect 8067 23613 8079 23647
rect 8021 23607 8079 23613
rect 6730 23536 6736 23588
rect 6788 23536 6794 23588
rect 8036 23576 8064 23607
rect 8478 23604 8484 23656
rect 8536 23644 8542 23656
rect 8536 23616 9674 23644
rect 8536 23604 8542 23616
rect 8665 23579 8723 23585
rect 8665 23576 8677 23579
rect 8036 23548 8677 23576
rect 8665 23545 8677 23548
rect 8711 23545 8723 23579
rect 8665 23539 8723 23545
rect 6362 23508 6368 23520
rect 6323 23480 6368 23508
rect 6362 23468 6368 23480
rect 6420 23468 6426 23520
rect 6914 23468 6920 23520
rect 6972 23508 6978 23520
rect 8110 23508 8116 23520
rect 6972 23480 8116 23508
rect 6972 23468 6978 23480
rect 8110 23468 8116 23480
rect 8168 23468 8174 23520
rect 9398 23508 9404 23520
rect 9359 23480 9404 23508
rect 9398 23468 9404 23480
rect 9456 23468 9462 23520
rect 9646 23508 9674 23616
rect 11716 23576 11744 23675
rect 11790 23656 11796 23708
rect 11848 23656 11854 23708
rect 11885 23681 11897 23715
rect 11931 23681 11943 23715
rect 11885 23675 11943 23681
rect 11900 23644 11928 23675
rect 11974 23672 11980 23724
rect 12032 23721 12038 23724
rect 12032 23715 12061 23721
rect 12049 23681 12061 23715
rect 12032 23675 12061 23681
rect 12032 23672 12038 23675
rect 12158 23672 12164 23724
rect 12216 23712 12222 23724
rect 12406 23712 12434 23752
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 15473 23783 15531 23789
rect 15473 23780 15485 23783
rect 14700 23752 15485 23780
rect 14700 23740 14706 23752
rect 15473 23749 15485 23752
rect 15519 23749 15531 23783
rect 16574 23780 16580 23792
rect 15473 23743 15531 23749
rect 15580 23752 16580 23780
rect 12805 23715 12863 23721
rect 12805 23712 12817 23715
rect 12216 23684 12261 23712
rect 12406 23684 12817 23712
rect 12216 23672 12222 23684
rect 12805 23681 12817 23684
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 12894 23672 12900 23724
rect 12952 23712 12958 23724
rect 13061 23715 13119 23721
rect 13061 23712 13073 23715
rect 12952 23684 13073 23712
rect 12952 23672 12958 23684
rect 13061 23681 13073 23684
rect 13107 23681 13119 23715
rect 13061 23675 13119 23681
rect 15286 23672 15292 23724
rect 15344 23721 15350 23724
rect 15580 23721 15608 23752
rect 16574 23740 16580 23752
rect 16632 23780 16638 23792
rect 17218 23780 17224 23792
rect 16632 23752 17224 23780
rect 16632 23740 16638 23752
rect 17218 23740 17224 23752
rect 17276 23740 17282 23792
rect 17310 23740 17316 23792
rect 17368 23780 17374 23792
rect 17862 23780 17868 23792
rect 17368 23752 17868 23780
rect 17368 23740 17374 23752
rect 17862 23740 17868 23752
rect 17920 23780 17926 23792
rect 26145 23783 26203 23789
rect 26145 23780 26157 23783
rect 17920 23752 21864 23780
rect 23322 23752 26157 23780
rect 17920 23740 17926 23752
rect 15344 23715 15366 23721
rect 15354 23681 15366 23715
rect 15344 23675 15366 23681
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23681 15623 23715
rect 16666 23712 16672 23724
rect 16627 23684 16672 23712
rect 15565 23675 15623 23681
rect 15344 23672 15350 23675
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 16850 23712 16856 23724
rect 16811 23684 16856 23712
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 18708 23721 18736 23752
rect 18426 23715 18484 23721
rect 18426 23712 18438 23715
rect 17696 23684 18438 23712
rect 16761 23647 16819 23653
rect 11900 23616 12011 23644
rect 11882 23576 11888 23588
rect 11716 23548 11888 23576
rect 11882 23536 11888 23548
rect 11940 23536 11946 23588
rect 10594 23508 10600 23520
rect 9646 23480 10600 23508
rect 10594 23468 10600 23480
rect 10652 23508 10658 23520
rect 11983 23508 12011 23616
rect 16761 23613 16773 23647
rect 16807 23644 16819 23647
rect 17696 23644 17724 23684
rect 18426 23681 18438 23684
rect 18472 23681 18484 23715
rect 18426 23675 18484 23681
rect 18693 23715 18751 23721
rect 18693 23681 18705 23715
rect 18739 23681 18751 23715
rect 18693 23675 18751 23681
rect 19242 23672 19248 23724
rect 19300 23712 19306 23724
rect 19613 23715 19671 23721
rect 19613 23712 19625 23715
rect 19300 23684 19625 23712
rect 19300 23672 19306 23684
rect 19613 23681 19625 23684
rect 19659 23681 19671 23715
rect 19613 23675 19671 23681
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23712 19855 23715
rect 19978 23712 19984 23724
rect 19843 23684 19984 23712
rect 19843 23681 19855 23684
rect 19797 23675 19855 23681
rect 19978 23672 19984 23684
rect 20036 23672 20042 23724
rect 20530 23712 20536 23724
rect 20491 23684 20536 23712
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 20622 23672 20628 23724
rect 20680 23712 20686 23724
rect 21836 23721 21864 23752
rect 26145 23749 26157 23752
rect 26191 23749 26203 23783
rect 26326 23780 26332 23792
rect 26145 23743 26203 23749
rect 26252 23752 26332 23780
rect 20717 23715 20775 23721
rect 20717 23712 20729 23715
rect 20680 23684 20729 23712
rect 20680 23672 20686 23684
rect 20717 23681 20729 23684
rect 20763 23681 20775 23715
rect 20717 23675 20775 23681
rect 21821 23715 21879 23721
rect 21821 23681 21833 23715
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 23382 23672 23388 23724
rect 23440 23712 23446 23724
rect 23842 23712 23848 23724
rect 23440 23684 23848 23712
rect 23440 23672 23446 23684
rect 23842 23672 23848 23684
rect 23900 23712 23906 23724
rect 24305 23715 24363 23721
rect 24305 23712 24317 23715
rect 23900 23684 24317 23712
rect 23900 23672 23906 23684
rect 24305 23681 24317 23684
rect 24351 23681 24363 23715
rect 24578 23712 24584 23724
rect 24539 23684 24584 23712
rect 24305 23675 24363 23681
rect 16807 23616 17724 23644
rect 16807 23613 16819 23616
rect 16761 23607 16819 23613
rect 20346 23604 20352 23656
rect 20404 23644 20410 23656
rect 20441 23647 20499 23653
rect 20441 23644 20453 23647
rect 20404 23616 20453 23644
rect 20404 23604 20410 23616
rect 20441 23613 20453 23616
rect 20487 23613 20499 23647
rect 20441 23607 20499 23613
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22152 23616 22197 23644
rect 22152 23604 22158 23616
rect 23658 23604 23664 23656
rect 23716 23604 23722 23656
rect 24320 23644 24348 23675
rect 24578 23672 24584 23684
rect 24636 23672 24642 23724
rect 24670 23672 24676 23724
rect 24728 23712 24734 23724
rect 26252 23721 26280 23752
rect 26326 23740 26332 23752
rect 26384 23780 26390 23792
rect 26384 23752 30788 23780
rect 26384 23740 26390 23752
rect 30760 23721 30788 23752
rect 25409 23715 25467 23721
rect 25409 23712 25421 23715
rect 24728 23684 25421 23712
rect 24728 23672 24734 23684
rect 25409 23681 25421 23684
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 26237 23715 26295 23721
rect 26237 23681 26249 23715
rect 26283 23681 26295 23715
rect 26237 23675 26295 23681
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23681 27491 23715
rect 27433 23675 27491 23681
rect 30745 23715 30803 23721
rect 30745 23681 30757 23715
rect 30791 23712 30803 23715
rect 31018 23712 31024 23724
rect 30791 23684 31024 23712
rect 30791 23681 30803 23684
rect 30745 23675 30803 23681
rect 25041 23647 25099 23653
rect 25041 23644 25053 23647
rect 24320 23616 25053 23644
rect 25041 23613 25053 23616
rect 25087 23613 25099 23647
rect 25590 23644 25596 23656
rect 25551 23616 25596 23644
rect 25041 23607 25099 23613
rect 25590 23604 25596 23616
rect 25648 23604 25654 23656
rect 12066 23536 12072 23588
rect 12124 23576 12130 23588
rect 12526 23576 12532 23588
rect 12124 23548 12532 23576
rect 12124 23536 12130 23548
rect 12526 23536 12532 23548
rect 12584 23536 12590 23588
rect 14090 23536 14096 23588
rect 14148 23576 14154 23588
rect 14185 23579 14243 23585
rect 14185 23576 14197 23579
rect 14148 23548 14197 23576
rect 14148 23536 14154 23548
rect 14185 23545 14197 23548
rect 14231 23545 14243 23579
rect 23676 23576 23704 23604
rect 27448 23576 27476 23675
rect 31018 23672 31024 23684
rect 31076 23672 31082 23724
rect 31726 23644 31754 23820
rect 32766 23808 32772 23820
rect 32824 23808 32830 23860
rect 34514 23848 34520 23860
rect 32876 23820 34520 23848
rect 32876 23721 32904 23820
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 34882 23808 34888 23860
rect 34940 23848 34946 23860
rect 37366 23848 37372 23860
rect 34940 23820 35572 23848
rect 37327 23820 37372 23848
rect 34940 23808 34946 23820
rect 34330 23780 34336 23792
rect 33980 23752 34336 23780
rect 32861 23715 32919 23721
rect 32861 23681 32873 23715
rect 32907 23681 32919 23715
rect 33502 23712 33508 23724
rect 33463 23684 33508 23712
rect 32861 23675 32919 23681
rect 33502 23672 33508 23684
rect 33560 23672 33566 23724
rect 33980 23721 34008 23752
rect 34330 23740 34336 23752
rect 34388 23740 34394 23792
rect 35544 23780 35572 23820
rect 37366 23808 37372 23820
rect 37424 23808 37430 23860
rect 35544 23752 37964 23780
rect 33965 23715 34023 23721
rect 33965 23681 33977 23715
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 35342 23672 35348 23724
rect 35400 23672 35406 23724
rect 36265 23715 36323 23721
rect 36265 23681 36277 23715
rect 36311 23681 36323 23715
rect 37274 23712 37280 23724
rect 37235 23684 37280 23712
rect 36265 23675 36323 23681
rect 23676 23548 27476 23576
rect 27540 23616 31754 23644
rect 14185 23539 14243 23545
rect 13170 23508 13176 23520
rect 10652 23480 13176 23508
rect 10652 23468 10658 23480
rect 13170 23468 13176 23480
rect 13228 23468 13234 23520
rect 17313 23511 17371 23517
rect 17313 23477 17325 23511
rect 17359 23508 17371 23511
rect 17494 23508 17500 23520
rect 17359 23480 17500 23508
rect 17359 23477 17371 23480
rect 17313 23471 17371 23477
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 20162 23468 20168 23520
rect 20220 23508 20226 23520
rect 23290 23508 23296 23520
rect 20220 23480 23296 23508
rect 20220 23468 20226 23480
rect 23290 23468 23296 23480
rect 23348 23508 23354 23520
rect 23569 23511 23627 23517
rect 23569 23508 23581 23511
rect 23348 23480 23581 23508
rect 23348 23468 23354 23480
rect 23569 23477 23581 23480
rect 23615 23477 23627 23511
rect 23569 23471 23627 23477
rect 23750 23468 23756 23520
rect 23808 23508 23814 23520
rect 27540 23508 27568 23616
rect 33686 23604 33692 23656
rect 33744 23644 33750 23656
rect 34241 23647 34299 23653
rect 34241 23644 34253 23647
rect 33744 23616 34253 23644
rect 33744 23604 33750 23616
rect 34241 23613 34253 23616
rect 34287 23613 34299 23647
rect 34241 23607 34299 23613
rect 34330 23604 34336 23656
rect 34388 23644 34394 23656
rect 36280 23644 36308 23675
rect 37274 23672 37280 23684
rect 37332 23672 37338 23724
rect 37936 23721 37964 23752
rect 37921 23715 37979 23721
rect 37921 23681 37933 23715
rect 37967 23681 37979 23715
rect 37921 23675 37979 23681
rect 37458 23644 37464 23656
rect 34388 23616 37464 23644
rect 34388 23604 34394 23616
rect 37458 23604 37464 23616
rect 37516 23604 37522 23656
rect 30929 23579 30987 23585
rect 30929 23545 30941 23579
rect 30975 23576 30987 23579
rect 31938 23576 31944 23588
rect 30975 23548 31944 23576
rect 30975 23545 30987 23548
rect 30929 23539 30987 23545
rect 31938 23536 31944 23548
rect 31996 23536 32002 23588
rect 36078 23576 36084 23588
rect 35544 23548 36084 23576
rect 23808 23480 27568 23508
rect 33413 23511 33471 23517
rect 23808 23468 23814 23480
rect 33413 23477 33425 23511
rect 33459 23508 33471 23511
rect 35544 23508 35572 23548
rect 36078 23536 36084 23548
rect 36136 23536 36142 23588
rect 35710 23508 35716 23520
rect 33459 23480 35572 23508
rect 35671 23480 35716 23508
rect 33459 23477 33471 23480
rect 33413 23471 33471 23477
rect 35710 23468 35716 23480
rect 35768 23468 35774 23520
rect 36354 23508 36360 23520
rect 36315 23480 36360 23508
rect 36354 23468 36360 23480
rect 36412 23468 36418 23520
rect 36538 23468 36544 23520
rect 36596 23508 36602 23520
rect 38013 23511 38071 23517
rect 38013 23508 38025 23511
rect 36596 23480 38025 23508
rect 36596 23468 36602 23480
rect 38013 23477 38025 23480
rect 38059 23477 38071 23511
rect 38013 23471 38071 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 6641 23307 6699 23313
rect 6641 23273 6653 23307
rect 6687 23304 6699 23307
rect 8846 23304 8852 23316
rect 6687 23276 8852 23304
rect 6687 23273 6699 23276
rect 6641 23267 6699 23273
rect 8846 23264 8852 23276
rect 8904 23304 8910 23316
rect 10321 23307 10379 23313
rect 8904 23276 10272 23304
rect 8904 23264 8910 23276
rect 7742 23168 7748 23180
rect 7703 23140 7748 23168
rect 7742 23128 7748 23140
rect 7800 23128 7806 23180
rect 10244 23168 10272 23276
rect 10321 23273 10333 23307
rect 10367 23304 10379 23307
rect 10410 23304 10416 23316
rect 10367 23276 10416 23304
rect 10367 23273 10379 23276
rect 10321 23267 10379 23273
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 11241 23307 11299 23313
rect 11241 23273 11253 23307
rect 11287 23304 11299 23307
rect 12342 23304 12348 23316
rect 11287 23276 12348 23304
rect 11287 23273 11299 23276
rect 11241 23267 11299 23273
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 12894 23304 12900 23316
rect 12855 23276 12900 23304
rect 12894 23264 12900 23276
rect 12952 23264 12958 23316
rect 15473 23307 15531 23313
rect 15473 23304 15485 23307
rect 15396 23276 15485 23304
rect 11149 23171 11207 23177
rect 10244 23140 10916 23168
rect 4338 23060 4344 23112
rect 4396 23100 4402 23112
rect 4614 23100 4620 23112
rect 4396 23072 4620 23100
rect 4396 23060 4402 23072
rect 4614 23060 4620 23072
rect 4672 23100 4678 23112
rect 5261 23103 5319 23109
rect 5261 23100 5273 23103
rect 4672 23072 5273 23100
rect 4672 23060 4678 23072
rect 5261 23069 5273 23072
rect 5307 23069 5319 23103
rect 5261 23063 5319 23069
rect 5528 23103 5586 23109
rect 5528 23069 5540 23103
rect 5574 23100 5586 23103
rect 6362 23100 6368 23112
rect 5574 23072 6368 23100
rect 5574 23069 5586 23072
rect 5528 23063 5586 23069
rect 6362 23060 6368 23072
rect 6420 23060 6426 23112
rect 7469 23103 7527 23109
rect 7469 23069 7481 23103
rect 7515 23100 7527 23103
rect 7834 23100 7840 23112
rect 7515 23072 7840 23100
rect 7515 23069 7527 23072
rect 7469 23063 7527 23069
rect 7834 23060 7840 23072
rect 7892 23060 7898 23112
rect 8938 23100 8944 23112
rect 8899 23072 8944 23100
rect 8938 23060 8944 23072
rect 8996 23060 9002 23112
rect 10410 23060 10416 23112
rect 10468 23100 10474 23112
rect 10781 23103 10839 23109
rect 10781 23100 10793 23103
rect 10468 23072 10793 23100
rect 10468 23060 10474 23072
rect 10781 23069 10793 23072
rect 10827 23069 10839 23103
rect 10888 23100 10916 23140
rect 11149 23137 11161 23171
rect 11195 23168 11207 23171
rect 11974 23168 11980 23180
rect 11195 23140 11980 23168
rect 11195 23137 11207 23140
rect 11149 23131 11207 23137
rect 11974 23128 11980 23140
rect 12032 23128 12038 23180
rect 14182 23168 14188 23180
rect 13096 23140 14188 23168
rect 11241 23103 11299 23109
rect 11241 23100 11253 23103
rect 10888 23072 11253 23100
rect 10781 23063 10839 23069
rect 11241 23069 11253 23072
rect 11287 23069 11299 23103
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 11241 23063 11299 23069
rect 11348 23072 12081 23100
rect 8754 22992 8760 23044
rect 8812 23032 8818 23044
rect 9186 23035 9244 23041
rect 9186 23032 9198 23035
rect 8812 23004 9198 23032
rect 8812 22992 8818 23004
rect 9186 23001 9198 23004
rect 9232 23001 9244 23035
rect 11348 23032 11376 23072
rect 12069 23069 12081 23072
rect 12115 23069 12127 23103
rect 12069 23063 12127 23069
rect 12161 23103 12219 23109
rect 12161 23069 12173 23103
rect 12207 23100 12219 23103
rect 12342 23100 12348 23112
rect 12207 23072 12348 23100
rect 12207 23069 12219 23072
rect 12161 23063 12219 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 13096 23109 13124 23140
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 15013 23171 15071 23177
rect 15013 23168 15025 23171
rect 14292 23140 15025 23168
rect 13081 23103 13139 23109
rect 13081 23069 13093 23103
rect 13127 23069 13139 23103
rect 13262 23100 13268 23112
rect 13223 23072 13268 23100
rect 13081 23063 13139 23069
rect 13262 23060 13268 23072
rect 13320 23060 13326 23112
rect 13354 23060 13360 23112
rect 13412 23109 13418 23112
rect 13412 23103 13441 23109
rect 13429 23069 13441 23103
rect 13412 23063 13441 23069
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23100 13599 23103
rect 13814 23100 13820 23112
rect 13587 23072 13820 23100
rect 13587 23069 13599 23072
rect 13541 23063 13599 23069
rect 13412 23060 13418 23063
rect 13814 23060 13820 23072
rect 13872 23100 13878 23112
rect 14090 23100 14096 23112
rect 13872 23072 14096 23100
rect 13872 23060 13878 23072
rect 14090 23060 14096 23072
rect 14148 23100 14154 23112
rect 14292 23100 14320 23140
rect 15013 23137 15025 23140
rect 15059 23168 15071 23171
rect 15396 23168 15424 23276
rect 15473 23273 15485 23276
rect 15519 23273 15531 23307
rect 16850 23304 16856 23316
rect 16811 23276 16856 23304
rect 15473 23267 15531 23273
rect 16850 23264 16856 23276
rect 16908 23264 16914 23316
rect 19058 23264 19064 23316
rect 19116 23304 19122 23316
rect 21450 23304 21456 23316
rect 19116 23276 21456 23304
rect 19116 23264 19122 23276
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 22005 23307 22063 23313
rect 22005 23273 22017 23307
rect 22051 23304 22063 23307
rect 22094 23304 22100 23316
rect 22051 23276 22100 23304
rect 22051 23273 22063 23276
rect 22005 23267 22063 23273
rect 22094 23264 22100 23276
rect 22152 23264 22158 23316
rect 34514 23264 34520 23316
rect 34572 23304 34578 23316
rect 35434 23304 35440 23316
rect 34572 23276 35440 23304
rect 34572 23264 34578 23276
rect 35434 23264 35440 23276
rect 35492 23264 35498 23316
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 19426 23236 19432 23248
rect 17092 23208 19432 23236
rect 17092 23196 17098 23208
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 21361 23239 21419 23245
rect 21361 23205 21373 23239
rect 21407 23236 21419 23239
rect 21407 23208 22324 23236
rect 21407 23205 21419 23208
rect 21361 23199 21419 23205
rect 15059 23140 15424 23168
rect 15059 23137 15071 23140
rect 15013 23131 15071 23137
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 15565 23171 15623 23177
rect 15565 23168 15577 23171
rect 15528 23140 15577 23168
rect 15528 23128 15534 23140
rect 15565 23137 15577 23140
rect 15611 23137 15623 23171
rect 15565 23131 15623 23137
rect 14642 23100 14648 23112
rect 14148 23072 14320 23100
rect 14603 23072 14648 23100
rect 14148 23060 14154 23072
rect 14642 23060 14648 23072
rect 14700 23060 14706 23112
rect 11882 23032 11888 23044
rect 9186 22995 9244 23001
rect 10796 23004 11376 23032
rect 11843 23004 11888 23032
rect 10796 22976 10824 23004
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 13170 23032 13176 23044
rect 13131 23004 13176 23032
rect 13170 22992 13176 23004
rect 13228 22992 13234 23044
rect 13998 23032 14004 23044
rect 13648 23004 14004 23032
rect 10778 22924 10784 22976
rect 10836 22924 10842 22976
rect 11422 22964 11428 22976
rect 11383 22936 11428 22964
rect 11422 22924 11428 22936
rect 11480 22924 11486 22976
rect 12158 22924 12164 22976
rect 12216 22964 12222 22976
rect 12253 22967 12311 22973
rect 12253 22964 12265 22967
rect 12216 22936 12265 22964
rect 12216 22924 12222 22936
rect 12253 22933 12265 22936
rect 12299 22933 12311 22967
rect 12253 22927 12311 22933
rect 12437 22967 12495 22973
rect 12437 22933 12449 22967
rect 12483 22964 12495 22967
rect 13648 22964 13676 23004
rect 13998 22992 14004 23004
rect 14056 23032 14062 23044
rect 14737 23035 14795 23041
rect 14737 23032 14749 23035
rect 14056 23004 14749 23032
rect 14056 22992 14062 23004
rect 14737 23001 14749 23004
rect 14783 23001 14795 23035
rect 15470 23032 15476 23044
rect 15431 23004 15476 23032
rect 14737 22995 14795 23001
rect 15470 22992 15476 23004
rect 15528 22992 15534 23044
rect 12483 22936 13676 22964
rect 14461 22967 14519 22973
rect 12483 22933 12495 22936
rect 12437 22927 12495 22933
rect 14461 22933 14473 22967
rect 14507 22964 14519 22967
rect 14550 22964 14556 22976
rect 14507 22936 14556 22964
rect 14507 22933 14519 22936
rect 14461 22927 14519 22933
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 14829 22967 14887 22973
rect 14829 22933 14841 22967
rect 14875 22964 14887 22967
rect 15580 22964 15608 23131
rect 16390 23128 16396 23180
rect 16448 23168 16454 23180
rect 19981 23171 20039 23177
rect 16448 23140 17448 23168
rect 16448 23128 16454 23140
rect 15746 23100 15752 23112
rect 15707 23072 15752 23100
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17034 23100 17040 23112
rect 16816 23072 17040 23100
rect 16816 23060 16822 23072
rect 17034 23060 17040 23072
rect 17092 23100 17098 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 17092 23072 17141 23100
rect 17092 23060 17098 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 17313 23103 17371 23109
rect 17313 23069 17325 23103
rect 17359 23097 17371 23103
rect 17420 23097 17448 23140
rect 19981 23137 19993 23171
rect 20027 23168 20039 23171
rect 20530 23168 20536 23180
rect 20027 23140 20536 23168
rect 20027 23137 20039 23140
rect 19981 23131 20039 23137
rect 20530 23128 20536 23140
rect 20588 23168 20594 23180
rect 22296 23177 22324 23208
rect 24578 23196 24584 23248
rect 24636 23236 24642 23248
rect 25590 23236 25596 23248
rect 24636 23208 25596 23236
rect 24636 23196 24642 23208
rect 25590 23196 25596 23208
rect 25648 23236 25654 23248
rect 25648 23208 29684 23236
rect 25648 23196 25654 23208
rect 22189 23171 22247 23177
rect 22189 23168 22201 23171
rect 20588 23140 22201 23168
rect 20588 23128 20594 23140
rect 22189 23137 22201 23140
rect 22235 23137 22247 23171
rect 22189 23131 22247 23137
rect 22281 23171 22339 23177
rect 22281 23137 22293 23171
rect 22327 23137 22339 23171
rect 22281 23131 22339 23137
rect 22373 23171 22431 23177
rect 22373 23137 22385 23171
rect 22419 23168 22431 23171
rect 23382 23168 23388 23180
rect 22419 23140 23388 23168
rect 22419 23137 22431 23140
rect 22373 23131 22431 23137
rect 23382 23128 23388 23140
rect 23440 23128 23446 23180
rect 26234 23168 26240 23180
rect 23584 23140 26240 23168
rect 17359 23069 17448 23097
rect 17313 23063 17371 23069
rect 17236 22976 17264 23063
rect 17494 23060 17500 23112
rect 17552 23100 17558 23112
rect 17954 23100 17960 23112
rect 17552 23072 17597 23100
rect 17915 23072 17960 23100
rect 17552 23060 17558 23072
rect 17954 23060 17960 23072
rect 18012 23060 18018 23112
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23100 18199 23103
rect 18230 23100 18236 23112
rect 18187 23072 18236 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 19426 23060 19432 23112
rect 19484 23100 19490 23112
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 19484 23072 19533 23100
rect 19484 23060 19490 23072
rect 19521 23069 19533 23072
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23100 19855 23103
rect 20070 23100 20076 23112
rect 19843 23072 20076 23100
rect 19843 23069 19855 23072
rect 19797 23063 19855 23069
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20625 23103 20683 23109
rect 20625 23100 20637 23103
rect 20220 23072 20637 23100
rect 20220 23060 20226 23072
rect 20625 23069 20637 23072
rect 20671 23069 20683 23103
rect 21174 23100 21180 23112
rect 21135 23072 21180 23100
rect 20625 23063 20683 23069
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 21269 23103 21327 23109
rect 21269 23069 21281 23103
rect 21315 23100 21327 23103
rect 21358 23100 21364 23112
rect 21315 23072 21364 23100
rect 21315 23069 21327 23072
rect 21269 23063 21327 23069
rect 21358 23060 21364 23072
rect 21416 23060 21422 23112
rect 21545 23103 21603 23109
rect 21545 23069 21557 23103
rect 21591 23100 21603 23103
rect 22465 23103 22523 23109
rect 21591 23072 22094 23100
rect 21591 23069 21603 23072
rect 21545 23063 21603 23069
rect 22066 23032 22094 23072
rect 22465 23069 22477 23103
rect 22511 23100 22523 23103
rect 23584 23100 23612 23140
rect 26234 23128 26240 23140
rect 26292 23128 26298 23180
rect 29546 23168 29552 23180
rect 26436 23140 27752 23168
rect 29507 23140 29552 23168
rect 22511 23072 23612 23100
rect 23661 23103 23719 23109
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 25038 23100 25044 23112
rect 23707 23072 25044 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 25406 23060 25412 23112
rect 25464 23100 25470 23112
rect 26436 23109 26464 23140
rect 25593 23103 25651 23109
rect 25593 23100 25605 23103
rect 25464 23072 25605 23100
rect 25464 23060 25470 23072
rect 25593 23069 25605 23072
rect 25639 23100 25651 23103
rect 26421 23103 26479 23109
rect 26421 23100 26433 23103
rect 25639 23072 26433 23100
rect 25639 23069 25651 23072
rect 25593 23063 25651 23069
rect 26421 23069 26433 23072
rect 26467 23069 26479 23103
rect 27062 23100 27068 23112
rect 27023 23072 27068 23100
rect 26421 23063 26479 23069
rect 27062 23060 27068 23072
rect 27120 23060 27126 23112
rect 27724 23109 27752 23140
rect 29546 23128 29552 23140
rect 29604 23128 29610 23180
rect 29656 23168 29684 23208
rect 30834 23196 30840 23248
rect 30892 23236 30898 23248
rect 30892 23208 32168 23236
rect 30892 23196 30898 23208
rect 32030 23168 32036 23180
rect 29656 23140 31754 23168
rect 31991 23140 32036 23168
rect 27709 23103 27767 23109
rect 27709 23069 27721 23103
rect 27755 23069 27767 23103
rect 27709 23063 27767 23069
rect 23382 23032 23388 23044
rect 22066 23004 23388 23032
rect 23382 22992 23388 23004
rect 23440 22992 23446 23044
rect 23845 23035 23903 23041
rect 23845 23001 23857 23035
rect 23891 23032 23903 23035
rect 24397 23035 24455 23041
rect 24397 23032 24409 23035
rect 23891 23004 24409 23032
rect 23891 23001 23903 23004
rect 23845 22995 23903 23001
rect 24397 23001 24409 23004
rect 24443 23001 24455 23035
rect 24578 23032 24584 23044
rect 24539 23004 24584 23032
rect 24397 22995 24455 23001
rect 24578 22992 24584 23004
rect 24636 22992 24642 23044
rect 24946 23032 24952 23044
rect 24907 23004 24952 23032
rect 24946 22992 24952 23004
rect 25004 22992 25010 23044
rect 25774 23032 25780 23044
rect 25056 23004 25780 23032
rect 14875 22936 15608 22964
rect 14875 22933 14887 22936
rect 14829 22927 14887 22933
rect 15654 22924 15660 22976
rect 15712 22964 15718 22976
rect 15933 22967 15991 22973
rect 15933 22964 15945 22967
rect 15712 22936 15945 22964
rect 15712 22924 15718 22936
rect 15933 22933 15945 22936
rect 15979 22933 15991 22967
rect 15933 22927 15991 22933
rect 17218 22924 17224 22976
rect 17276 22924 17282 22976
rect 18046 22964 18052 22976
rect 18007 22936 18052 22964
rect 18046 22924 18052 22936
rect 18104 22924 18110 22976
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 19613 22967 19671 22973
rect 19613 22964 19625 22967
rect 18932 22936 19625 22964
rect 18932 22924 18938 22936
rect 19613 22933 19625 22936
rect 19659 22933 19671 22967
rect 19613 22927 19671 22933
rect 20438 22924 20444 22976
rect 20496 22964 20502 22976
rect 20533 22967 20591 22973
rect 20533 22964 20545 22967
rect 20496 22936 20545 22964
rect 20496 22924 20502 22936
rect 20533 22933 20545 22936
rect 20579 22933 20591 22967
rect 20533 22927 20591 22933
rect 23477 22967 23535 22973
rect 23477 22933 23489 22967
rect 23523 22964 23535 22967
rect 24302 22964 24308 22976
rect 23523 22936 24308 22964
rect 23523 22933 23535 22936
rect 23477 22927 23535 22933
rect 24302 22924 24308 22936
rect 24360 22924 24366 22976
rect 24486 22924 24492 22976
rect 24544 22964 24550 22976
rect 24673 22967 24731 22973
rect 24673 22964 24685 22967
rect 24544 22936 24685 22964
rect 24544 22924 24550 22936
rect 24673 22933 24685 22936
rect 24719 22933 24731 22967
rect 24673 22927 24731 22933
rect 24765 22967 24823 22973
rect 24765 22933 24777 22967
rect 24811 22964 24823 22967
rect 25056 22964 25084 23004
rect 25774 22992 25780 23004
rect 25832 22992 25838 23044
rect 29454 22992 29460 23044
rect 29512 23032 29518 23044
rect 29825 23035 29883 23041
rect 29825 23032 29837 23035
rect 29512 23004 29837 23032
rect 29512 22992 29518 23004
rect 29825 23001 29837 23004
rect 29871 23001 29883 23035
rect 29825 22995 29883 23001
rect 30374 22992 30380 23044
rect 30432 22992 30438 23044
rect 31726 23032 31754 23140
rect 32030 23128 32036 23140
rect 32088 23128 32094 23180
rect 32140 23168 32168 23208
rect 36354 23168 36360 23180
rect 32140 23140 35296 23168
rect 36315 23140 36360 23168
rect 33410 23060 33416 23112
rect 33468 23060 33474 23112
rect 35268 23109 35296 23140
rect 36354 23128 36360 23140
rect 36412 23128 36418 23180
rect 38010 23168 38016 23180
rect 37971 23140 38016 23168
rect 38010 23128 38016 23140
rect 38068 23128 38074 23180
rect 35253 23103 35311 23109
rect 35253 23069 35265 23103
rect 35299 23069 35311 23103
rect 35253 23063 35311 23069
rect 31846 23032 31852 23044
rect 31726 23004 31852 23032
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 32306 23032 32312 23044
rect 32267 23004 32312 23032
rect 32306 22992 32312 23004
rect 32364 22992 32370 23044
rect 25498 22964 25504 22976
rect 24811 22936 25084 22964
rect 25459 22936 25504 22964
rect 24811 22933 24823 22936
rect 24765 22927 24823 22933
rect 25498 22924 25504 22936
rect 25556 22924 25562 22976
rect 26510 22964 26516 22976
rect 26471 22936 26516 22964
rect 26510 22924 26516 22936
rect 26568 22924 26574 22976
rect 27246 22964 27252 22976
rect 27207 22936 27252 22964
rect 27246 22924 27252 22936
rect 27304 22924 27310 22976
rect 27798 22964 27804 22976
rect 27759 22936 27804 22964
rect 27798 22924 27804 22936
rect 27856 22924 27862 22976
rect 31294 22964 31300 22976
rect 31255 22936 31300 22964
rect 31294 22924 31300 22936
rect 31352 22924 31358 22976
rect 33042 22924 33048 22976
rect 33100 22964 33106 22976
rect 33781 22967 33839 22973
rect 33781 22964 33793 22967
rect 33100 22936 33793 22964
rect 33100 22924 33106 22936
rect 33781 22933 33793 22936
rect 33827 22933 33839 22967
rect 35268 22964 35296 23063
rect 35986 23060 35992 23112
rect 36044 23100 36050 23112
rect 36173 23103 36231 23109
rect 36173 23100 36185 23103
rect 36044 23072 36185 23100
rect 36044 23060 36050 23072
rect 36173 23069 36185 23072
rect 36219 23069 36231 23103
rect 36173 23063 36231 23069
rect 36170 22964 36176 22976
rect 35268 22936 36176 22964
rect 33781 22927 33839 22933
rect 36170 22924 36176 22936
rect 36228 22924 36234 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 8754 22760 8760 22772
rect 8715 22732 8760 22760
rect 8754 22720 8760 22732
rect 8812 22720 8818 22772
rect 9398 22720 9404 22772
rect 9456 22760 9462 22772
rect 9493 22763 9551 22769
rect 9493 22760 9505 22763
rect 9456 22732 9505 22760
rect 9456 22720 9462 22732
rect 9493 22729 9505 22732
rect 9539 22729 9551 22763
rect 9493 22723 9551 22729
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 10597 22763 10655 22769
rect 10597 22760 10609 22763
rect 9732 22732 10609 22760
rect 9732 22720 9738 22732
rect 10597 22729 10609 22732
rect 10643 22729 10655 22763
rect 11885 22763 11943 22769
rect 11885 22760 11897 22763
rect 10597 22723 10655 22729
rect 11348 22732 11897 22760
rect 6733 22695 6791 22701
rect 6733 22661 6745 22695
rect 6779 22692 6791 22695
rect 7561 22695 7619 22701
rect 7561 22692 7573 22695
rect 6779 22664 7573 22692
rect 6779 22661 6791 22664
rect 6733 22655 6791 22661
rect 7561 22661 7573 22664
rect 7607 22661 7619 22695
rect 7561 22655 7619 22661
rect 7834 22652 7840 22704
rect 7892 22692 7898 22704
rect 9585 22695 9643 22701
rect 9585 22692 9597 22695
rect 7892 22664 9597 22692
rect 7892 22652 7898 22664
rect 9585 22661 9597 22664
rect 9631 22661 9643 22695
rect 9585 22655 9643 22661
rect 9769 22695 9827 22701
rect 9769 22661 9781 22695
rect 9815 22692 9827 22695
rect 11348 22692 11376 22732
rect 11885 22729 11897 22732
rect 11931 22760 11943 22763
rect 11974 22760 11980 22772
rect 11931 22732 11980 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12069 22763 12127 22769
rect 12069 22729 12081 22763
rect 12115 22760 12127 22763
rect 12250 22760 12256 22772
rect 12115 22732 12256 22760
rect 12115 22729 12127 22732
rect 12069 22723 12127 22729
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 12526 22760 12532 22772
rect 12487 22732 12532 22760
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 13170 22720 13176 22772
rect 13228 22760 13234 22772
rect 13541 22763 13599 22769
rect 13541 22760 13553 22763
rect 13228 22732 13553 22760
rect 13228 22720 13234 22732
rect 13541 22729 13553 22732
rect 13587 22729 13599 22763
rect 13541 22723 13599 22729
rect 16942 22720 16948 22772
rect 17000 22760 17006 22772
rect 17129 22763 17187 22769
rect 17129 22760 17141 22763
rect 17000 22732 17141 22760
rect 17000 22720 17006 22732
rect 17129 22729 17141 22732
rect 17175 22729 17187 22763
rect 17129 22723 17187 22729
rect 18969 22763 19027 22769
rect 18969 22729 18981 22763
rect 19015 22760 19027 22763
rect 19613 22763 19671 22769
rect 19613 22760 19625 22763
rect 19015 22732 19625 22760
rect 19015 22729 19027 22732
rect 18969 22723 19027 22729
rect 19613 22729 19625 22732
rect 19659 22760 19671 22763
rect 19659 22732 19932 22760
rect 19659 22729 19671 22732
rect 19613 22723 19671 22729
rect 19904 22704 19932 22732
rect 24302 22720 24308 22772
rect 24360 22760 24366 22772
rect 29454 22760 29460 22772
rect 24360 22732 26188 22760
rect 29415 22732 29460 22760
rect 24360 22720 24366 22732
rect 9815 22664 11376 22692
rect 9815 22661 9827 22664
rect 9769 22655 9827 22661
rect 11422 22652 11428 22704
rect 11480 22692 11486 22704
rect 11480 22664 13584 22692
rect 11480 22652 11486 22664
rect 4338 22624 4344 22636
rect 4299 22596 4344 22624
rect 4338 22584 4344 22596
rect 4396 22584 4402 22636
rect 4608 22627 4666 22633
rect 4608 22593 4620 22627
rect 4654 22624 4666 22627
rect 6365 22627 6423 22633
rect 6365 22624 6377 22627
rect 4654 22596 6377 22624
rect 4654 22593 4666 22596
rect 4608 22587 4666 22593
rect 6365 22593 6377 22596
rect 6411 22593 6423 22627
rect 6546 22624 6552 22636
rect 6507 22596 6552 22624
rect 6365 22587 6423 22593
rect 6546 22584 6552 22596
rect 6604 22584 6610 22636
rect 6638 22584 6644 22636
rect 6696 22624 6702 22636
rect 6696 22596 6789 22624
rect 6696 22584 6702 22596
rect 6822 22584 6828 22636
rect 6880 22633 6886 22636
rect 6880 22627 6909 22633
rect 6897 22624 6909 22627
rect 7653 22627 7711 22633
rect 6897 22596 7604 22624
rect 6897 22593 6909 22596
rect 6880 22587 6909 22593
rect 6880 22584 6886 22587
rect 6656 22488 6684 22584
rect 7006 22556 7012 22568
rect 6967 22528 7012 22556
rect 7006 22516 7012 22528
rect 7064 22516 7070 22568
rect 7576 22556 7604 22596
rect 7653 22593 7665 22627
rect 7699 22624 7711 22627
rect 7742 22624 7748 22636
rect 7699 22596 7748 22624
rect 7699 22593 7711 22596
rect 7653 22587 7711 22593
rect 7742 22584 7748 22596
rect 7800 22584 7806 22636
rect 8205 22627 8263 22633
rect 8205 22593 8217 22627
rect 8251 22624 8263 22627
rect 8294 22624 8300 22636
rect 8251 22596 8300 22624
rect 8251 22593 8263 22596
rect 8205 22587 8263 22593
rect 8294 22584 8300 22596
rect 8352 22584 8358 22636
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22593 8539 22627
rect 8481 22587 8539 22593
rect 8386 22556 8392 22568
rect 7576 22528 8392 22556
rect 8386 22516 8392 22528
rect 8444 22556 8450 22568
rect 8496 22556 8524 22587
rect 8570 22584 8576 22636
rect 8628 22624 8634 22636
rect 9401 22627 9459 22633
rect 9401 22624 9413 22627
rect 8628 22596 8673 22624
rect 8864 22596 9413 22624
rect 8628 22584 8634 22596
rect 8444 22528 8524 22556
rect 8444 22516 8450 22528
rect 7558 22488 7564 22500
rect 6656 22460 7564 22488
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 8478 22448 8484 22500
rect 8536 22488 8542 22500
rect 8864 22488 8892 22596
rect 9401 22593 9413 22596
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 10413 22627 10471 22633
rect 10413 22624 10425 22627
rect 10192 22596 10425 22624
rect 10192 22584 10198 22596
rect 10413 22593 10425 22596
rect 10459 22593 10471 22627
rect 10413 22587 10471 22593
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 10704 22556 10732 22587
rect 10778 22584 10784 22636
rect 10836 22624 10842 22636
rect 11701 22627 11759 22633
rect 10836 22596 10881 22624
rect 10836 22584 10842 22596
rect 11701 22593 11713 22627
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 12158 22624 12164 22636
rect 11839 22596 12164 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 11238 22556 11244 22568
rect 10704 22528 11244 22556
rect 11238 22516 11244 22528
rect 11296 22556 11302 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11296 22528 11529 22556
rect 11296 22516 11302 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 11716 22556 11744 22587
rect 12158 22584 12164 22596
rect 12216 22624 12222 22636
rect 12989 22627 13047 22633
rect 12989 22624 13001 22627
rect 12216 22596 13001 22624
rect 12216 22584 12222 22596
rect 12989 22593 13001 22596
rect 13035 22593 13047 22627
rect 12989 22587 13047 22593
rect 12710 22556 12716 22568
rect 11716 22528 11816 22556
rect 12671 22528 12716 22556
rect 11517 22519 11575 22525
rect 8536 22460 8892 22488
rect 9217 22491 9275 22497
rect 8536 22448 8542 22460
rect 9217 22457 9229 22491
rect 9263 22457 9275 22491
rect 9217 22451 9275 22457
rect 5721 22423 5779 22429
rect 5721 22389 5733 22423
rect 5767 22420 5779 22423
rect 5902 22420 5908 22432
rect 5767 22392 5908 22420
rect 5767 22389 5779 22392
rect 5721 22383 5779 22389
rect 5902 22380 5908 22392
rect 5960 22380 5966 22432
rect 8294 22420 8300 22432
rect 8255 22392 8300 22420
rect 8294 22380 8300 22392
rect 8352 22380 8358 22432
rect 8846 22380 8852 22432
rect 8904 22420 8910 22432
rect 9232 22420 9260 22451
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 11146 22488 11152 22500
rect 10468 22460 11152 22488
rect 10468 22448 10474 22460
rect 11146 22448 11152 22460
rect 11204 22488 11210 22500
rect 11788 22488 11816 22528
rect 12710 22516 12716 22528
rect 12768 22516 12774 22568
rect 12805 22559 12863 22565
rect 12805 22525 12817 22559
rect 12851 22525 12863 22559
rect 12805 22519 12863 22525
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22525 12955 22559
rect 13556 22556 13584 22664
rect 13630 22652 13636 22704
rect 13688 22692 13694 22704
rect 13909 22695 13967 22701
rect 13909 22692 13921 22695
rect 13688 22664 13921 22692
rect 13688 22652 13694 22664
rect 13909 22661 13921 22664
rect 13955 22661 13967 22695
rect 14458 22692 14464 22704
rect 14419 22664 14464 22692
rect 13909 22655 13967 22661
rect 14458 22652 14464 22664
rect 14516 22652 14522 22704
rect 15746 22652 15752 22704
rect 15804 22692 15810 22704
rect 16206 22692 16212 22704
rect 15804 22664 16212 22692
rect 15804 22652 15810 22664
rect 16206 22652 16212 22664
rect 16264 22692 16270 22704
rect 17494 22692 17500 22704
rect 16264 22664 17500 22692
rect 16264 22652 16270 22664
rect 13725 22627 13783 22633
rect 13725 22593 13737 22627
rect 13771 22624 13783 22627
rect 13814 22624 13820 22636
rect 13771 22596 13820 22624
rect 13771 22593 13783 22596
rect 13725 22587 13783 22593
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 13998 22624 14004 22636
rect 13959 22596 14004 22624
rect 13998 22584 14004 22596
rect 14056 22584 14062 22636
rect 14366 22584 14372 22636
rect 14424 22624 14430 22636
rect 14645 22627 14703 22633
rect 14645 22624 14657 22627
rect 14424 22596 14657 22624
rect 14424 22584 14430 22596
rect 14645 22593 14657 22596
rect 14691 22593 14703 22627
rect 15381 22627 15439 22633
rect 15381 22624 15393 22627
rect 14645 22587 14703 22593
rect 14752 22596 15393 22624
rect 14752 22556 14780 22596
rect 15381 22593 15393 22596
rect 15427 22593 15439 22627
rect 15654 22624 15660 22636
rect 15615 22596 15660 22624
rect 15381 22587 15439 22593
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 15838 22624 15844 22636
rect 15799 22596 15844 22624
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 16114 22624 16120 22636
rect 16075 22596 16120 22624
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 16960 22633 16988 22664
rect 17494 22652 17500 22664
rect 17552 22652 17558 22704
rect 18874 22692 18880 22704
rect 18835 22664 18880 22692
rect 18874 22652 18880 22664
rect 18932 22652 18938 22704
rect 19886 22652 19892 22704
rect 19944 22652 19950 22704
rect 22738 22692 22744 22704
rect 20824 22664 22744 22692
rect 16945 22627 17003 22633
rect 16945 22593 16957 22627
rect 16991 22593 17003 22627
rect 17218 22624 17224 22636
rect 17179 22596 17224 22624
rect 16945 22587 17003 22593
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 18138 22624 18144 22636
rect 18099 22596 18144 22624
rect 18138 22584 18144 22596
rect 18196 22584 18202 22636
rect 20824 22633 20852 22664
rect 22738 22652 22744 22664
rect 22796 22652 22802 22704
rect 25498 22692 25504 22704
rect 25254 22664 25504 22692
rect 25498 22652 25504 22664
rect 25556 22652 25562 22704
rect 18693 22627 18751 22633
rect 18693 22593 18705 22627
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 18969 22627 19027 22633
rect 18969 22593 18981 22627
rect 19015 22624 19027 22627
rect 20809 22627 20867 22633
rect 20809 22624 20821 22627
rect 19015 22596 20821 22624
rect 19015 22593 19027 22596
rect 18969 22587 19027 22593
rect 20809 22593 20821 22596
rect 20855 22593 20867 22627
rect 20809 22587 20867 22593
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22624 21143 22627
rect 21358 22624 21364 22636
rect 21131 22596 21364 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 13556 22528 14780 22556
rect 15289 22559 15347 22565
rect 12897 22519 12955 22525
rect 15289 22525 15301 22559
rect 15335 22556 15347 22559
rect 18708 22556 18736 22587
rect 21358 22584 21364 22596
rect 21416 22584 21422 22636
rect 26160 22633 26188 22732
rect 29454 22720 29460 22732
rect 29512 22720 29518 22772
rect 33410 22720 33416 22772
rect 33468 22760 33474 22772
rect 33505 22763 33563 22769
rect 33505 22760 33517 22763
rect 33468 22732 33517 22760
rect 33468 22720 33474 22732
rect 33505 22729 33517 22732
rect 33551 22729 33563 22763
rect 33505 22723 33563 22729
rect 27246 22692 27252 22704
rect 27207 22664 27252 22692
rect 27246 22652 27252 22664
rect 27304 22652 27310 22704
rect 27798 22652 27804 22704
rect 27856 22652 27862 22704
rect 28552 22664 37320 22692
rect 26145 22627 26203 22633
rect 26145 22593 26157 22627
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 19426 22556 19432 22568
rect 15335 22528 19432 22556
rect 15335 22525 15347 22528
rect 15289 22519 15347 22525
rect 12820 22488 12848 22519
rect 11204 22460 12848 22488
rect 11204 22448 11210 22460
rect 10686 22420 10692 22432
rect 8904 22392 9260 22420
rect 10647 22392 10692 22420
rect 8904 22380 8910 22392
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 12342 22380 12348 22432
rect 12400 22420 12406 22432
rect 12912 22420 12940 22519
rect 19426 22516 19432 22528
rect 19484 22516 19490 22568
rect 19978 22556 19984 22568
rect 19939 22528 19984 22556
rect 19978 22516 19984 22528
rect 20036 22556 20042 22568
rect 22278 22556 22284 22568
rect 20036 22528 22284 22556
rect 20036 22516 20042 22528
rect 22278 22516 22284 22528
rect 22336 22556 22342 22568
rect 22465 22559 22523 22565
rect 22465 22556 22477 22559
rect 22336 22528 22477 22556
rect 22336 22516 22342 22528
rect 22465 22525 22477 22528
rect 22511 22525 22523 22559
rect 22465 22519 22523 22525
rect 22741 22559 22799 22565
rect 22741 22525 22753 22559
rect 22787 22525 22799 22559
rect 22741 22519 22799 22525
rect 16666 22448 16672 22500
rect 16724 22488 16730 22500
rect 16945 22491 17003 22497
rect 16945 22488 16957 22491
rect 16724 22460 16957 22488
rect 16724 22448 16730 22460
rect 16945 22457 16957 22460
rect 16991 22457 17003 22491
rect 16945 22451 17003 22457
rect 20809 22491 20867 22497
rect 20809 22457 20821 22491
rect 20855 22488 20867 22491
rect 22554 22488 22560 22500
rect 20855 22460 22560 22488
rect 20855 22457 20867 22460
rect 20809 22451 20867 22457
rect 22554 22448 22560 22460
rect 22612 22448 22618 22500
rect 22646 22448 22652 22500
rect 22704 22488 22710 22500
rect 22756 22488 22784 22519
rect 23198 22516 23204 22568
rect 23256 22556 23262 22568
rect 23566 22556 23572 22568
rect 23256 22528 23572 22556
rect 23256 22516 23262 22528
rect 23566 22516 23572 22528
rect 23624 22556 23630 22568
rect 23753 22559 23811 22565
rect 23753 22556 23765 22559
rect 23624 22528 23765 22556
rect 23624 22516 23630 22528
rect 23753 22525 23765 22528
rect 23799 22525 23811 22559
rect 23753 22519 23811 22525
rect 24029 22559 24087 22565
rect 24029 22525 24041 22559
rect 24075 22556 24087 22559
rect 26973 22559 27031 22565
rect 26973 22556 26985 22559
rect 24075 22528 26004 22556
rect 24075 22525 24087 22528
rect 24029 22519 24087 22525
rect 23658 22488 23664 22500
rect 22704 22460 23664 22488
rect 22704 22448 22710 22460
rect 23658 22448 23664 22460
rect 23716 22448 23722 22500
rect 25976 22497 26004 22528
rect 26160 22528 26985 22556
rect 26160 22500 26188 22528
rect 26973 22525 26985 22528
rect 27019 22525 27031 22559
rect 26973 22519 27031 22525
rect 25961 22491 26019 22497
rect 25056 22460 25636 22488
rect 12400 22392 12940 22420
rect 12400 22380 12406 22392
rect 15286 22380 15292 22432
rect 15344 22420 15350 22432
rect 18049 22423 18107 22429
rect 18049 22420 18061 22423
rect 15344 22392 18061 22420
rect 15344 22380 15350 22392
rect 18049 22389 18061 22392
rect 18095 22389 18107 22423
rect 18049 22383 18107 22389
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19429 22423 19487 22429
rect 19429 22420 19441 22423
rect 19392 22392 19441 22420
rect 19392 22380 19398 22392
rect 19429 22389 19441 22392
rect 19475 22389 19487 22423
rect 19429 22383 19487 22389
rect 19610 22380 19616 22432
rect 19668 22420 19674 22432
rect 21174 22420 21180 22432
rect 19668 22392 21180 22420
rect 19668 22380 19674 22392
rect 21174 22380 21180 22392
rect 21232 22380 21238 22432
rect 23014 22380 23020 22432
rect 23072 22420 23078 22432
rect 25056 22420 25084 22460
rect 25498 22420 25504 22432
rect 23072 22392 25084 22420
rect 25459 22392 25504 22420
rect 23072 22380 23078 22392
rect 25498 22380 25504 22392
rect 25556 22380 25562 22432
rect 25608 22420 25636 22460
rect 25961 22457 25973 22491
rect 26007 22457 26019 22491
rect 25961 22451 26019 22457
rect 26142 22448 26148 22500
rect 26200 22448 26206 22500
rect 28552 22420 28580 22664
rect 29270 22624 29276 22636
rect 29231 22596 29276 22624
rect 29270 22584 29276 22596
rect 29328 22584 29334 22636
rect 30098 22624 30104 22636
rect 30059 22596 30104 22624
rect 30098 22584 30104 22596
rect 30156 22584 30162 22636
rect 30466 22584 30472 22636
rect 30524 22624 30530 22636
rect 30561 22627 30619 22633
rect 30561 22624 30573 22627
rect 30524 22596 30573 22624
rect 30524 22584 30530 22596
rect 30561 22593 30573 22596
rect 30607 22624 30619 22627
rect 30834 22624 30840 22636
rect 30607 22596 30840 22624
rect 30607 22593 30619 22596
rect 30561 22587 30619 22593
rect 30834 22584 30840 22596
rect 30892 22584 30898 22636
rect 32309 22627 32367 22633
rect 32309 22624 32321 22627
rect 31726 22596 32321 22624
rect 25608 22392 28580 22420
rect 28721 22423 28779 22429
rect 28721 22389 28733 22423
rect 28767 22420 28779 22423
rect 28994 22420 29000 22432
rect 28767 22392 29000 22420
rect 28767 22389 28779 22392
rect 28721 22383 28779 22389
rect 28994 22380 29000 22392
rect 29052 22380 29058 22432
rect 30006 22420 30012 22432
rect 29967 22392 30012 22420
rect 30006 22380 30012 22392
rect 30064 22380 30070 22432
rect 30098 22380 30104 22432
rect 30156 22420 30162 22432
rect 30745 22423 30803 22429
rect 30745 22420 30757 22423
rect 30156 22392 30757 22420
rect 30156 22380 30162 22392
rect 30745 22389 30757 22392
rect 30791 22420 30803 22423
rect 31726 22420 31754 22596
rect 32309 22593 32321 22596
rect 32355 22624 32367 22627
rect 32953 22627 33011 22633
rect 32953 22624 32965 22627
rect 32355 22596 32965 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 32953 22593 32965 22596
rect 32999 22624 33011 22627
rect 33413 22627 33471 22633
rect 33413 22624 33425 22627
rect 32999 22596 33425 22624
rect 32999 22593 33011 22596
rect 32953 22587 33011 22593
rect 33413 22593 33425 22596
rect 33459 22593 33471 22627
rect 33413 22587 33471 22593
rect 34425 22627 34483 22633
rect 34425 22593 34437 22627
rect 34471 22593 34483 22627
rect 34425 22587 34483 22593
rect 33870 22516 33876 22568
rect 33928 22556 33934 22568
rect 34149 22559 34207 22565
rect 34149 22556 34161 22559
rect 33928 22528 34161 22556
rect 33928 22516 33934 22528
rect 34149 22525 34161 22528
rect 34195 22525 34207 22559
rect 34149 22519 34207 22525
rect 31938 22448 31944 22500
rect 31996 22488 32002 22500
rect 32861 22491 32919 22497
rect 32861 22488 32873 22491
rect 31996 22460 32873 22488
rect 31996 22448 32002 22460
rect 32861 22457 32873 22460
rect 32907 22457 32919 22491
rect 32861 22451 32919 22457
rect 33778 22448 33784 22500
rect 33836 22488 33842 22500
rect 34333 22491 34391 22497
rect 34333 22488 34345 22491
rect 33836 22460 34345 22488
rect 33836 22448 33842 22460
rect 34333 22457 34345 22460
rect 34379 22457 34391 22491
rect 34440 22488 34468 22587
rect 34606 22584 34612 22636
rect 34664 22624 34670 22636
rect 37292 22633 37320 22664
rect 34885 22627 34943 22633
rect 34885 22624 34897 22627
rect 34664 22596 34897 22624
rect 34664 22584 34670 22596
rect 34885 22593 34897 22596
rect 34931 22593 34943 22627
rect 34885 22587 34943 22593
rect 37277 22627 37335 22633
rect 37277 22593 37289 22627
rect 37323 22593 37335 22627
rect 37277 22587 37335 22593
rect 37458 22584 37464 22636
rect 37516 22624 37522 22636
rect 37921 22627 37979 22633
rect 37921 22624 37933 22627
rect 37516 22596 37933 22624
rect 37516 22584 37522 22596
rect 37921 22593 37933 22596
rect 37967 22593 37979 22627
rect 37921 22587 37979 22593
rect 35069 22559 35127 22565
rect 35069 22525 35081 22559
rect 35115 22556 35127 22559
rect 36538 22556 36544 22568
rect 35115 22528 36544 22556
rect 35115 22525 35127 22528
rect 35069 22519 35127 22525
rect 36538 22516 36544 22528
rect 36596 22516 36602 22568
rect 36722 22556 36728 22568
rect 36683 22528 36728 22556
rect 36722 22516 36728 22528
rect 36780 22516 36786 22568
rect 36998 22516 37004 22568
rect 37056 22556 37062 22568
rect 37476 22556 37504 22584
rect 37056 22528 37504 22556
rect 37056 22516 37062 22528
rect 34440 22460 36400 22488
rect 34333 22451 34391 22457
rect 30791 22392 31754 22420
rect 30791 22389 30803 22392
rect 30745 22383 30803 22389
rect 32122 22380 32128 22432
rect 32180 22420 32186 22432
rect 32217 22423 32275 22429
rect 32217 22420 32229 22423
rect 32180 22392 32229 22420
rect 32180 22380 32186 22392
rect 32217 22389 32229 22392
rect 32263 22389 32275 22423
rect 32217 22383 32275 22389
rect 34425 22423 34483 22429
rect 34425 22389 34437 22423
rect 34471 22420 34483 22423
rect 34698 22420 34704 22432
rect 34471 22392 34704 22420
rect 34471 22389 34483 22392
rect 34425 22383 34483 22389
rect 34698 22380 34704 22392
rect 34756 22380 34762 22432
rect 36372 22420 36400 22460
rect 36446 22448 36452 22500
rect 36504 22488 36510 22500
rect 38013 22491 38071 22497
rect 38013 22488 38025 22491
rect 36504 22460 38025 22488
rect 36504 22448 36510 22460
rect 38013 22457 38025 22460
rect 38059 22457 38071 22491
rect 38013 22451 38071 22457
rect 37274 22420 37280 22432
rect 36372 22392 37280 22420
rect 37274 22380 37280 22392
rect 37332 22380 37338 22432
rect 37369 22423 37427 22429
rect 37369 22389 37381 22423
rect 37415 22420 37427 22423
rect 37918 22420 37924 22432
rect 37415 22392 37924 22420
rect 37415 22389 37427 22392
rect 37369 22383 37427 22389
rect 37918 22380 37924 22392
rect 37976 22380 37982 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 6641 22219 6699 22225
rect 6641 22185 6653 22219
rect 6687 22216 6699 22219
rect 7098 22216 7104 22228
rect 6687 22188 7104 22216
rect 6687 22185 6699 22188
rect 6641 22179 6699 22185
rect 7098 22176 7104 22188
rect 7156 22216 7162 22228
rect 7156 22188 7788 22216
rect 7156 22176 7162 22188
rect 7469 22151 7527 22157
rect 7469 22117 7481 22151
rect 7515 22148 7527 22151
rect 7650 22148 7656 22160
rect 7515 22120 7656 22148
rect 7515 22117 7527 22120
rect 7469 22111 7527 22117
rect 7650 22108 7656 22120
rect 7708 22108 7714 22160
rect 7760 22148 7788 22188
rect 8294 22176 8300 22228
rect 8352 22216 8358 22228
rect 9125 22219 9183 22225
rect 9125 22216 9137 22219
rect 8352 22188 9137 22216
rect 8352 22176 8358 22188
rect 9125 22185 9137 22188
rect 9171 22185 9183 22219
rect 10410 22216 10416 22228
rect 10371 22188 10416 22216
rect 9125 22179 9183 22185
rect 10410 22176 10416 22188
rect 10468 22176 10474 22228
rect 10594 22176 10600 22228
rect 10652 22176 10658 22228
rect 10686 22176 10692 22228
rect 10744 22216 10750 22228
rect 14182 22216 14188 22228
rect 10744 22188 14188 22216
rect 10744 22176 10750 22188
rect 14182 22176 14188 22188
rect 14240 22176 14246 22228
rect 14642 22176 14648 22228
rect 14700 22216 14706 22228
rect 15381 22219 15439 22225
rect 15381 22216 15393 22219
rect 14700 22188 15393 22216
rect 14700 22176 14706 22188
rect 15381 22185 15393 22188
rect 15427 22185 15439 22219
rect 15381 22179 15439 22185
rect 17681 22219 17739 22225
rect 17681 22185 17693 22219
rect 17727 22216 17739 22219
rect 17954 22216 17960 22228
rect 17727 22188 17960 22216
rect 17727 22185 17739 22188
rect 17681 22179 17739 22185
rect 17954 22176 17960 22188
rect 18012 22176 18018 22228
rect 20441 22219 20499 22225
rect 20441 22185 20453 22219
rect 20487 22216 20499 22219
rect 20530 22216 20536 22228
rect 20487 22188 20536 22216
rect 20487 22185 20499 22188
rect 20441 22179 20499 22185
rect 20530 22176 20536 22188
rect 20588 22176 20594 22228
rect 25038 22216 25044 22228
rect 24999 22188 25044 22216
rect 25038 22176 25044 22188
rect 25096 22176 25102 22228
rect 33042 22216 33048 22228
rect 28966 22188 31984 22216
rect 33003 22188 33048 22216
rect 7760 22120 7880 22148
rect 5902 22040 5908 22092
rect 5960 22080 5966 22092
rect 5960 22052 6868 22080
rect 5960 22040 5966 22052
rect 6362 22012 6368 22024
rect 6323 21984 6368 22012
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 6641 22015 6699 22021
rect 6641 21981 6653 22015
rect 6687 22012 6699 22015
rect 6730 22012 6736 22024
rect 6687 21984 6736 22012
rect 6687 21981 6699 21984
rect 6641 21975 6699 21981
rect 6730 21972 6736 21984
rect 6788 21972 6794 22024
rect 6840 22012 6868 22052
rect 7006 22012 7012 22024
rect 6840 21984 7012 22012
rect 7006 21972 7012 21984
rect 7064 22012 7070 22024
rect 7852 22021 7880 22120
rect 10612 22080 10640 22176
rect 11195 22151 11253 22157
rect 11195 22117 11207 22151
rect 11241 22148 11253 22151
rect 11330 22148 11336 22160
rect 11241 22120 11336 22148
rect 11241 22117 11253 22120
rect 11195 22111 11253 22117
rect 11330 22108 11336 22120
rect 11388 22108 11394 22160
rect 11974 22108 11980 22160
rect 12032 22148 12038 22160
rect 12032 22120 12940 22148
rect 12032 22108 12038 22120
rect 10686 22080 10692 22092
rect 10612 22052 10692 22080
rect 10686 22040 10692 22052
rect 10744 22040 10750 22092
rect 11256 22052 11836 22080
rect 11256 22024 11284 22052
rect 7653 22015 7711 22021
rect 7653 22012 7665 22015
rect 7064 21984 7665 22012
rect 7064 21972 7070 21984
rect 7653 21981 7665 21984
rect 7699 21981 7711 22015
rect 7653 21975 7711 21981
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8110 21972 8116 22024
rect 8168 22012 8174 22024
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8168 21984 8953 22012
rect 8168 21972 8174 21984
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 10226 22012 10232 22024
rect 9171 21984 10232 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10597 22015 10655 22021
rect 10597 21981 10609 22015
rect 10643 22012 10655 22015
rect 10778 22012 10784 22024
rect 10643 21984 10784 22012
rect 10643 21981 10655 21984
rect 10597 21975 10655 21981
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 11057 22015 11115 22021
rect 11057 21981 11069 22015
rect 11103 22012 11115 22015
rect 11238 22012 11244 22024
rect 11103 21984 11244 22012
rect 11103 21981 11115 21984
rect 11057 21975 11115 21981
rect 11238 21972 11244 21984
rect 11296 21972 11302 22024
rect 11330 21972 11336 22024
rect 11388 22012 11394 22024
rect 11514 22012 11520 22024
rect 11388 21984 11433 22012
rect 11475 21984 11520 22012
rect 11388 21972 11394 21984
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 11808 22012 11836 22052
rect 11882 22040 11888 22092
rect 11940 22080 11946 22092
rect 12253 22083 12311 22089
rect 12253 22080 12265 22083
rect 11940 22052 12265 22080
rect 11940 22040 11946 22052
rect 12253 22049 12265 22052
rect 12299 22049 12311 22083
rect 12912 22080 12940 22120
rect 14458 22108 14464 22160
rect 14516 22148 14522 22160
rect 16390 22148 16396 22160
rect 14516 22120 16396 22148
rect 14516 22108 14522 22120
rect 16390 22108 16396 22120
rect 16448 22148 16454 22160
rect 19610 22148 19616 22160
rect 16448 22120 16528 22148
rect 16448 22108 16454 22120
rect 13078 22080 13084 22092
rect 12912 22052 13084 22080
rect 12253 22043 12311 22049
rect 13078 22040 13084 22052
rect 13136 22080 13142 22092
rect 14093 22083 14151 22089
rect 14093 22080 14105 22083
rect 13136 22052 14105 22080
rect 13136 22040 13142 22052
rect 14093 22049 14105 22052
rect 14139 22049 14151 22083
rect 15746 22080 15752 22092
rect 15707 22052 15752 22080
rect 14093 22043 14151 22049
rect 15746 22040 15752 22052
rect 15804 22040 15810 22092
rect 12342 22012 12348 22024
rect 11808 21984 12348 22012
rect 12342 21972 12348 21984
rect 12400 22012 12406 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12400 21984 12541 22012
rect 12400 21972 12406 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 13630 21972 13636 22024
rect 13688 22012 13694 22024
rect 14369 22015 14427 22021
rect 14369 22012 14381 22015
rect 13688 21984 14381 22012
rect 13688 21972 13694 21984
rect 14369 21981 14381 21984
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 15470 21972 15476 22024
rect 15528 22012 15534 22024
rect 16500 22021 16528 22120
rect 19260 22120 19616 22148
rect 16945 22083 17003 22089
rect 16592 22052 16896 22080
rect 16592 22021 16620 22052
rect 15565 22015 15623 22021
rect 15565 22012 15577 22015
rect 15528 21984 15577 22012
rect 15528 21972 15534 21984
rect 15565 21981 15577 21984
rect 15611 21981 15623 22015
rect 15565 21975 15623 21981
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 16577 22015 16635 22021
rect 16577 21981 16589 22015
rect 16623 21981 16635 22015
rect 16577 21975 16635 21981
rect 8021 21947 8079 21953
rect 6840 21916 7972 21944
rect 6840 21885 6868 21916
rect 6825 21879 6883 21885
rect 6825 21845 6837 21879
rect 6871 21845 6883 21879
rect 7742 21876 7748 21888
rect 7703 21848 7748 21876
rect 6825 21839 6883 21845
rect 7742 21836 7748 21848
rect 7800 21836 7806 21888
rect 7944 21876 7972 21916
rect 8021 21913 8033 21947
rect 8067 21944 8079 21947
rect 8754 21944 8760 21956
rect 8067 21916 8760 21944
rect 8067 21913 8079 21916
rect 8021 21907 8079 21913
rect 8754 21904 8760 21916
rect 8812 21904 8818 21956
rect 15838 21944 15844 21956
rect 9600 21916 15844 21944
rect 9600 21876 9628 21916
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 16316 21944 16344 21975
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 16868 22012 16896 22052
rect 16945 22049 16957 22083
rect 16991 22080 17003 22083
rect 18230 22080 18236 22092
rect 16991 22052 18236 22080
rect 16991 22049 17003 22052
rect 16945 22043 17003 22049
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 17126 22012 17132 22024
rect 16724 21984 16769 22012
rect 16868 21984 17132 22012
rect 16724 21972 16730 21984
rect 17126 21972 17132 21984
rect 17184 22012 17190 22024
rect 17405 22015 17463 22021
rect 17405 22012 17417 22015
rect 17184 21984 17417 22012
rect 17184 21972 17190 21984
rect 17405 21981 17417 21984
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 22012 18659 22015
rect 19150 22012 19156 22024
rect 18647 21984 19156 22012
rect 18647 21981 18659 21984
rect 18601 21975 18659 21981
rect 19150 21972 19156 21984
rect 19208 21972 19214 22024
rect 19260 22021 19288 22120
rect 19610 22108 19616 22120
rect 19668 22108 19674 22160
rect 23566 22108 23572 22160
rect 23624 22108 23630 22160
rect 19886 22080 19892 22092
rect 19847 22052 19892 22080
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 20257 22083 20315 22089
rect 20257 22049 20269 22083
rect 20303 22080 20315 22083
rect 21358 22080 21364 22092
rect 20303 22052 21364 22080
rect 20303 22049 20315 22052
rect 20257 22043 20315 22049
rect 21358 22040 21364 22052
rect 21416 22080 21422 22092
rect 22005 22083 22063 22089
rect 22005 22080 22017 22083
rect 21416 22052 22017 22080
rect 21416 22040 21422 22052
rect 22005 22049 22017 22052
rect 22051 22080 22063 22083
rect 23584 22080 23612 22108
rect 25777 22083 25835 22089
rect 25777 22080 25789 22083
rect 22051 22052 23244 22080
rect 23584 22052 25789 22080
rect 22051 22049 22063 22052
rect 22005 22043 22063 22049
rect 19245 22015 19303 22021
rect 19245 21981 19257 22015
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 22278 22012 22284 22024
rect 22191 21984 22284 22012
rect 19429 21975 19487 21981
rect 16390 21944 16396 21956
rect 16303 21916 16396 21944
rect 16390 21904 16396 21916
rect 16448 21944 16454 21956
rect 17681 21947 17739 21953
rect 17681 21944 17693 21947
rect 16448 21916 17693 21944
rect 16448 21904 16454 21916
rect 17681 21913 17693 21916
rect 17727 21913 17739 21947
rect 18414 21944 18420 21956
rect 18375 21916 18420 21944
rect 17681 21907 17739 21913
rect 18414 21904 18420 21916
rect 18472 21904 18478 21956
rect 19444 21888 19472 21975
rect 22278 21972 22284 21984
rect 22336 22012 22342 22024
rect 22925 22015 22983 22021
rect 22925 22012 22937 22015
rect 22336 21984 22937 22012
rect 22336 21972 22342 21984
rect 22925 21981 22937 21984
rect 22971 21981 22983 22015
rect 22925 21975 22983 21981
rect 22738 21944 22744 21956
rect 22699 21916 22744 21944
rect 22738 21904 22744 21916
rect 22796 21904 22802 21956
rect 23014 21904 23020 21956
rect 23072 21944 23078 21956
rect 23109 21947 23167 21953
rect 23109 21944 23121 21947
rect 23072 21916 23121 21944
rect 23072 21904 23078 21916
rect 23109 21913 23121 21916
rect 23155 21913 23167 21947
rect 23216 21944 23244 22052
rect 25777 22049 25789 22052
rect 25823 22080 25835 22083
rect 26142 22080 26148 22092
rect 25823 22052 26148 22080
rect 25823 22049 25835 22052
rect 25777 22043 25835 22049
rect 26142 22040 26148 22052
rect 26200 22040 26206 22092
rect 27525 22083 27583 22089
rect 27525 22049 27537 22083
rect 27571 22080 27583 22083
rect 27706 22080 27712 22092
rect 27571 22052 27712 22080
rect 27571 22049 27583 22052
rect 27525 22043 27583 22049
rect 27706 22040 27712 22052
rect 27764 22040 27770 22092
rect 28966 22080 28994 22188
rect 29546 22108 29552 22160
rect 29604 22148 29610 22160
rect 31956 22148 31984 22188
rect 33042 22176 33048 22188
rect 33100 22176 33106 22228
rect 33778 22216 33784 22228
rect 33739 22188 33784 22216
rect 33778 22176 33784 22188
rect 33836 22176 33842 22228
rect 33965 22219 34023 22225
rect 33965 22185 33977 22219
rect 34011 22185 34023 22219
rect 33965 22179 34023 22185
rect 35345 22219 35403 22225
rect 35345 22185 35357 22219
rect 35391 22216 35403 22219
rect 35710 22216 35716 22228
rect 35391 22188 35716 22216
rect 35391 22185 35403 22188
rect 35345 22179 35403 22185
rect 33980 22148 34008 22179
rect 35710 22176 35716 22188
rect 35768 22176 35774 22228
rect 35986 22176 35992 22228
rect 36044 22216 36050 22228
rect 37182 22216 37188 22228
rect 36044 22188 37188 22216
rect 36044 22176 36050 22188
rect 37182 22176 37188 22188
rect 37240 22176 37246 22228
rect 35434 22148 35440 22160
rect 29604 22120 30328 22148
rect 31956 22120 35440 22148
rect 29604 22108 29610 22120
rect 28184 22052 28994 22080
rect 30300 22080 30328 22120
rect 35434 22108 35440 22120
rect 35492 22108 35498 22160
rect 30469 22083 30527 22089
rect 30469 22080 30481 22083
rect 30300 22052 30481 22080
rect 23290 21972 23296 22024
rect 23348 22012 23354 22024
rect 23569 22015 23627 22021
rect 23569 22012 23581 22015
rect 23348 21984 23581 22012
rect 23348 21972 23354 21984
rect 23569 21981 23581 21984
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 23658 21972 23664 22024
rect 23716 22012 23722 22024
rect 23753 22015 23811 22021
rect 23753 22012 23765 22015
rect 23716 21984 23765 22012
rect 23716 21972 23722 21984
rect 23753 21981 23765 21984
rect 23799 21981 23811 22015
rect 23753 21975 23811 21981
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 22012 24915 22015
rect 25498 22012 25504 22024
rect 24903 21984 25504 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 24780 21944 24808 21975
rect 25498 21972 25504 21984
rect 25556 21972 25562 22024
rect 27982 21972 27988 22024
rect 28040 22012 28046 22024
rect 28184 22021 28212 22052
rect 30469 22049 30481 22052
rect 30515 22049 30527 22083
rect 30469 22043 30527 22049
rect 31110 22040 31116 22092
rect 31168 22080 31174 22092
rect 32861 22083 32919 22089
rect 32861 22080 32873 22083
rect 31168 22052 32873 22080
rect 31168 22040 31174 22052
rect 32861 22049 32873 22052
rect 32907 22049 32919 22083
rect 35894 22080 35900 22092
rect 32861 22043 32919 22049
rect 33060 22052 35900 22080
rect 28169 22015 28227 22021
rect 28169 22012 28181 22015
rect 28040 21984 28181 22012
rect 28040 21972 28046 21984
rect 28169 21981 28181 21984
rect 28215 21981 28227 22015
rect 28350 22012 28356 22024
rect 28311 21984 28356 22012
rect 28169 21975 28227 21981
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 28997 22015 29055 22021
rect 28997 21981 29009 22015
rect 29043 22012 29055 22015
rect 29086 22012 29092 22024
rect 29043 21984 29092 22012
rect 29043 21981 29055 21984
rect 28997 21975 29055 21981
rect 29086 21972 29092 21984
rect 29144 21972 29150 22024
rect 30009 22015 30067 22021
rect 30009 21981 30021 22015
rect 30055 22012 30067 22015
rect 30098 22012 30104 22024
rect 30055 21984 30104 22012
rect 30055 21981 30067 21984
rect 30009 21975 30067 21981
rect 30098 21972 30104 21984
rect 30156 21972 30162 22024
rect 33060 22021 33088 22052
rect 35894 22040 35900 22052
rect 35952 22040 35958 22092
rect 37458 22080 37464 22092
rect 37419 22052 37464 22080
rect 37458 22040 37464 22052
rect 37516 22040 37522 22092
rect 37918 22080 37924 22092
rect 37879 22052 37924 22080
rect 37918 22040 37924 22052
rect 37976 22040 37982 22092
rect 38105 22083 38163 22089
rect 38105 22049 38117 22083
rect 38151 22080 38163 22083
rect 38194 22080 38200 22092
rect 38151 22052 38200 22080
rect 38151 22049 38163 22052
rect 38105 22043 38163 22049
rect 38194 22040 38200 22052
rect 38252 22040 38258 22092
rect 33045 22015 33103 22021
rect 33045 21981 33057 22015
rect 33091 21981 33103 22015
rect 33045 21975 33103 21981
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 35069 22015 35127 22021
rect 35069 22012 35081 22015
rect 34848 21984 35081 22012
rect 34848 21972 34854 21984
rect 35069 21981 35081 21984
rect 35115 21981 35127 22015
rect 35069 21975 35127 21981
rect 35161 22015 35219 22021
rect 35161 21981 35173 22015
rect 35207 22012 35219 22015
rect 35207 21984 35756 22012
rect 35207 21981 35219 21984
rect 35161 21975 35219 21981
rect 24946 21944 24952 21956
rect 23216 21916 24952 21944
rect 23109 21907 23167 21913
rect 24946 21904 24952 21916
rect 25004 21904 25010 21956
rect 26053 21947 26111 21953
rect 26053 21913 26065 21947
rect 26099 21944 26111 21947
rect 26326 21944 26332 21956
rect 26099 21916 26332 21944
rect 26099 21913 26111 21916
rect 26053 21907 26111 21913
rect 26326 21904 26332 21916
rect 26384 21904 26390 21956
rect 26510 21904 26516 21956
rect 26568 21904 26574 21956
rect 29917 21947 29975 21953
rect 29917 21913 29929 21947
rect 29963 21944 29975 21947
rect 30374 21944 30380 21956
rect 29963 21916 30380 21944
rect 29963 21913 29975 21916
rect 29917 21907 29975 21913
rect 30374 21904 30380 21916
rect 30432 21904 30438 21956
rect 30742 21944 30748 21956
rect 30703 21916 30748 21944
rect 30742 21904 30748 21916
rect 30800 21904 30806 21956
rect 32122 21944 32128 21956
rect 31970 21916 32128 21944
rect 32122 21904 32128 21916
rect 32180 21904 32186 21956
rect 32769 21947 32827 21953
rect 32769 21913 32781 21947
rect 32815 21913 32827 21947
rect 32769 21907 32827 21913
rect 34149 21947 34207 21953
rect 34149 21913 34161 21947
rect 34195 21944 34207 21947
rect 35176 21944 35204 21975
rect 35342 21944 35348 21956
rect 34195 21916 35204 21944
rect 35303 21916 35348 21944
rect 34195 21913 34207 21916
rect 34149 21907 34207 21913
rect 7944 21848 9628 21876
rect 11517 21879 11575 21885
rect 11517 21845 11529 21879
rect 11563 21876 11575 21879
rect 11606 21876 11612 21888
rect 11563 21848 11612 21876
rect 11563 21845 11575 21848
rect 11517 21839 11575 21845
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 14826 21836 14832 21888
rect 14884 21876 14890 21888
rect 17497 21879 17555 21885
rect 17497 21876 17509 21879
rect 14884 21848 17509 21876
rect 14884 21836 14890 21848
rect 17497 21845 17509 21848
rect 17543 21845 17555 21879
rect 19242 21876 19248 21888
rect 19203 21848 19248 21876
rect 17497 21839 17555 21845
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 19426 21836 19432 21888
rect 19484 21836 19490 21888
rect 20070 21876 20076 21888
rect 20031 21848 20076 21876
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 23753 21879 23811 21885
rect 23753 21845 23765 21879
rect 23799 21876 23811 21879
rect 23842 21876 23848 21888
rect 23799 21848 23848 21876
rect 23799 21845 23811 21848
rect 23753 21839 23811 21845
rect 23842 21836 23848 21848
rect 23900 21836 23906 21888
rect 24394 21876 24400 21888
rect 24355 21848 24400 21876
rect 24394 21836 24400 21848
rect 24452 21836 24458 21888
rect 24578 21836 24584 21888
rect 24636 21876 24642 21888
rect 26234 21876 26240 21888
rect 24636 21848 26240 21876
rect 24636 21836 24642 21848
rect 26234 21836 26240 21848
rect 26292 21836 26298 21888
rect 27614 21836 27620 21888
rect 27672 21876 27678 21888
rect 28169 21879 28227 21885
rect 28169 21876 28181 21879
rect 27672 21848 28181 21876
rect 27672 21836 27678 21848
rect 28169 21845 28181 21848
rect 28215 21845 28227 21879
rect 28902 21876 28908 21888
rect 28863 21848 28908 21876
rect 28169 21839 28227 21845
rect 28902 21836 28908 21848
rect 28960 21836 28966 21888
rect 32214 21876 32220 21888
rect 32175 21848 32220 21876
rect 32214 21836 32220 21848
rect 32272 21876 32278 21888
rect 32784 21876 32812 21907
rect 35342 21904 35348 21916
rect 35400 21904 35406 21956
rect 35728 21944 35756 21984
rect 37274 21944 37280 21956
rect 35728 21916 37280 21944
rect 37274 21904 37280 21916
rect 37332 21904 37338 21956
rect 33226 21876 33232 21888
rect 32272 21848 32812 21876
rect 33187 21848 33232 21876
rect 32272 21836 32278 21848
rect 33226 21836 33232 21848
rect 33284 21836 33290 21888
rect 33962 21885 33968 21888
rect 33949 21879 33968 21885
rect 33949 21845 33961 21879
rect 33949 21839 33968 21845
rect 33962 21836 33968 21839
rect 34020 21836 34026 21888
rect 34054 21836 34060 21888
rect 34112 21876 34118 21888
rect 34885 21879 34943 21885
rect 34885 21876 34897 21879
rect 34112 21848 34897 21876
rect 34112 21836 34118 21848
rect 34885 21845 34897 21848
rect 34931 21845 34943 21879
rect 34885 21839 34943 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 4614 21632 4620 21684
rect 4672 21632 4678 21684
rect 5721 21675 5779 21681
rect 5721 21641 5733 21675
rect 5767 21672 5779 21675
rect 6362 21672 6368 21684
rect 5767 21644 6368 21672
rect 5767 21641 5779 21644
rect 5721 21635 5779 21641
rect 6362 21632 6368 21644
rect 6420 21632 6426 21684
rect 7558 21632 7564 21684
rect 7616 21672 7622 21684
rect 10505 21675 10563 21681
rect 7616 21644 8892 21672
rect 7616 21632 7622 21644
rect 4632 21604 4660 21632
rect 7944 21613 7972 21644
rect 7653 21607 7711 21613
rect 7653 21604 7665 21607
rect 4356 21576 4660 21604
rect 6104 21576 7665 21604
rect 4356 21545 4384 21576
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21505 4399 21539
rect 4341 21499 4399 21505
rect 4608 21539 4666 21545
rect 4608 21505 4620 21539
rect 4654 21536 4666 21539
rect 6104 21536 6132 21576
rect 7653 21573 7665 21576
rect 7699 21573 7711 21607
rect 7653 21567 7711 21573
rect 7929 21607 7987 21613
rect 7929 21573 7941 21607
rect 7975 21573 7987 21607
rect 7929 21567 7987 21573
rect 8018 21564 8024 21616
rect 8076 21604 8082 21616
rect 8159 21607 8217 21613
rect 8076 21576 8121 21604
rect 8076 21564 8082 21576
rect 8159 21573 8171 21607
rect 8205 21604 8217 21607
rect 8386 21604 8392 21616
rect 8205 21576 8392 21604
rect 8205 21573 8217 21576
rect 8159 21567 8217 21573
rect 8386 21564 8392 21576
rect 8444 21564 8450 21616
rect 6362 21536 6368 21548
rect 4654 21508 6132 21536
rect 6323 21508 6368 21536
rect 4654 21505 4666 21508
rect 4608 21499 4666 21505
rect 6362 21496 6368 21508
rect 6420 21496 6426 21548
rect 7834 21536 7840 21548
rect 7795 21508 7840 21536
rect 7834 21496 7840 21508
rect 7892 21496 7898 21548
rect 6638 21468 6644 21480
rect 6599 21440 6644 21468
rect 6638 21428 6644 21440
rect 6696 21468 6702 21480
rect 7742 21468 7748 21480
rect 6696 21440 7748 21468
rect 6696 21428 6702 21440
rect 7742 21428 7748 21440
rect 7800 21468 7806 21480
rect 8297 21471 8355 21477
rect 8297 21468 8309 21471
rect 7800 21440 8309 21468
rect 7800 21428 7806 21440
rect 8297 21437 8309 21440
rect 8343 21437 8355 21471
rect 8297 21431 8355 21437
rect 5442 21360 5448 21412
rect 5500 21400 5506 21412
rect 8018 21400 8024 21412
rect 5500 21372 8024 21400
rect 5500 21360 5506 21372
rect 8018 21360 8024 21372
rect 8076 21360 8082 21412
rect 6730 21292 6736 21344
rect 6788 21332 6794 21344
rect 8754 21332 8760 21344
rect 6788 21304 8760 21332
rect 6788 21292 6794 21304
rect 8754 21292 8760 21304
rect 8812 21292 8818 21344
rect 8864 21332 8892 21644
rect 10505 21641 10517 21675
rect 10551 21672 10563 21675
rect 10778 21672 10784 21684
rect 10551 21644 10784 21672
rect 10551 21641 10563 21644
rect 10505 21635 10563 21641
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 12897 21675 12955 21681
rect 12897 21672 12909 21675
rect 11940 21644 12909 21672
rect 11940 21632 11946 21644
rect 12897 21641 12909 21644
rect 12943 21641 12955 21675
rect 12897 21635 12955 21641
rect 13998 21632 14004 21684
rect 14056 21672 14062 21684
rect 20254 21672 20260 21684
rect 14056 21644 20260 21672
rect 14056 21632 14062 21644
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 23569 21675 23627 21681
rect 23569 21641 23581 21675
rect 23615 21672 23627 21675
rect 30466 21672 30472 21684
rect 23615 21644 24624 21672
rect 23615 21641 23627 21644
rect 23569 21635 23627 21641
rect 17804 21607 17862 21613
rect 9140 21576 11560 21604
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9140 21477 9168 21576
rect 9392 21539 9450 21545
rect 9392 21505 9404 21539
rect 9438 21536 9450 21539
rect 10502 21536 10508 21548
rect 9438 21508 10508 21536
rect 9438 21505 9450 21508
rect 9392 21499 9450 21505
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 11532 21545 11560 21576
rect 17804 21573 17816 21607
rect 17850 21604 17862 21607
rect 18046 21604 18052 21616
rect 17850 21576 18052 21604
rect 17850 21573 17862 21576
rect 17804 21567 17862 21573
rect 18046 21564 18052 21576
rect 18104 21564 18110 21616
rect 18138 21564 18144 21616
rect 18196 21604 18202 21616
rect 18693 21607 18751 21613
rect 18693 21604 18705 21607
rect 18196 21576 18705 21604
rect 18196 21564 18202 21576
rect 18693 21573 18705 21576
rect 18739 21604 18751 21607
rect 19242 21604 19248 21616
rect 18739 21576 19248 21604
rect 18739 21573 18751 21576
rect 18693 21567 18751 21573
rect 19242 21564 19248 21576
rect 19300 21564 19306 21616
rect 19613 21607 19671 21613
rect 19613 21573 19625 21607
rect 19659 21604 19671 21607
rect 20898 21604 20904 21616
rect 19659 21576 20904 21604
rect 19659 21573 19671 21576
rect 19613 21567 19671 21573
rect 20898 21564 20904 21576
rect 20956 21604 20962 21616
rect 24394 21604 24400 21616
rect 20956 21576 24400 21604
rect 20956 21564 20962 21576
rect 24394 21564 24400 21576
rect 24452 21564 24458 21616
rect 11517 21539 11575 21545
rect 11517 21505 11529 21539
rect 11563 21505 11575 21539
rect 11517 21499 11575 21505
rect 11606 21496 11612 21548
rect 11664 21536 11670 21548
rect 11773 21539 11831 21545
rect 11773 21536 11785 21539
rect 11664 21508 11785 21536
rect 11664 21496 11670 21508
rect 11773 21505 11785 21508
rect 11819 21505 11831 21539
rect 11773 21499 11831 21505
rect 12802 21496 12808 21548
rect 12860 21536 12866 21548
rect 13541 21539 13599 21545
rect 13541 21536 13553 21539
rect 12860 21508 13553 21536
rect 12860 21496 12866 21508
rect 13541 21505 13553 21508
rect 13587 21536 13599 21539
rect 13630 21536 13636 21548
rect 13587 21508 13636 21536
rect 13587 21505 13599 21508
rect 13541 21499 13599 21505
rect 13630 21496 13636 21508
rect 13688 21496 13694 21548
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21505 13783 21539
rect 13725 21499 13783 21505
rect 13909 21539 13967 21545
rect 13909 21505 13921 21539
rect 13955 21536 13967 21539
rect 14090 21536 14096 21548
rect 13955 21508 14096 21536
rect 13955 21505 13967 21508
rect 13909 21499 13967 21505
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 8996 21440 9137 21468
rect 8996 21428 9002 21440
rect 9125 21437 9137 21440
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 13170 21428 13176 21480
rect 13228 21468 13234 21480
rect 13740 21468 13768 21499
rect 14090 21496 14096 21508
rect 14148 21536 14154 21548
rect 14369 21539 14427 21545
rect 14369 21536 14381 21539
rect 14148 21508 14381 21536
rect 14148 21496 14154 21508
rect 14369 21505 14381 21508
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 15562 21536 15568 21548
rect 14599 21508 15568 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 15562 21496 15568 21508
rect 15620 21496 15626 21548
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 15933 21539 15991 21545
rect 15933 21536 15945 21539
rect 15896 21508 15945 21536
rect 15896 21496 15902 21508
rect 15933 21505 15945 21508
rect 15979 21505 15991 21539
rect 19334 21536 19340 21548
rect 19295 21508 19340 21536
rect 15933 21499 15991 21505
rect 19334 21496 19340 21508
rect 19392 21496 19398 21548
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21505 19487 21539
rect 19429 21499 19487 21505
rect 15102 21468 15108 21480
rect 13228 21440 15108 21468
rect 13228 21428 13234 21440
rect 14568 21412 14596 21440
rect 15102 21428 15108 21440
rect 15160 21428 15166 21480
rect 15749 21471 15807 21477
rect 15749 21437 15761 21471
rect 15795 21468 15807 21471
rect 16390 21468 16396 21480
rect 15795 21440 16396 21468
rect 15795 21437 15807 21440
rect 15749 21431 15807 21437
rect 16390 21428 16396 21440
rect 16448 21428 16454 21480
rect 18046 21468 18052 21480
rect 18007 21440 18052 21468
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 18598 21428 18604 21480
rect 18656 21468 18662 21480
rect 19058 21468 19064 21480
rect 18656 21440 19064 21468
rect 18656 21428 18662 21440
rect 19058 21428 19064 21440
rect 19116 21468 19122 21480
rect 19444 21468 19472 21499
rect 19978 21496 19984 21548
rect 20036 21536 20042 21548
rect 20257 21539 20315 21545
rect 20257 21536 20269 21539
rect 20036 21508 20269 21536
rect 20036 21496 20042 21508
rect 20257 21505 20269 21508
rect 20303 21505 20315 21539
rect 20438 21536 20444 21548
rect 20399 21508 20444 21536
rect 20257 21499 20315 21505
rect 20438 21496 20444 21508
rect 20496 21536 20502 21548
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20496 21508 21097 21536
rect 20496 21496 20502 21508
rect 21085 21505 21097 21508
rect 21131 21536 21143 21539
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21131 21508 21833 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 22097 21539 22155 21545
rect 22097 21505 22109 21539
rect 22143 21536 22155 21539
rect 22738 21536 22744 21548
rect 22143 21508 22744 21536
rect 22143 21505 22155 21508
rect 22097 21499 22155 21505
rect 22738 21496 22744 21508
rect 22796 21496 22802 21548
rect 23106 21496 23112 21548
rect 23164 21536 23170 21548
rect 24596 21545 24624 21644
rect 25608 21644 30472 21672
rect 24762 21564 24768 21616
rect 24820 21604 24826 21616
rect 25227 21607 25285 21613
rect 25227 21604 25239 21607
rect 24820 21576 25239 21604
rect 24820 21564 24826 21576
rect 25227 21573 25239 21576
rect 25273 21604 25285 21607
rect 25608 21604 25636 21644
rect 30466 21632 30472 21644
rect 30524 21632 30530 21684
rect 30745 21675 30803 21681
rect 30745 21641 30757 21675
rect 30791 21672 30803 21675
rect 30834 21672 30840 21684
rect 30791 21644 30840 21672
rect 30791 21641 30803 21644
rect 30745 21635 30803 21641
rect 30834 21632 30840 21644
rect 30892 21672 30898 21684
rect 31294 21672 31300 21684
rect 30892 21644 31300 21672
rect 30892 21632 30898 21644
rect 31294 21632 31300 21644
rect 31352 21632 31358 21684
rect 34514 21672 34520 21684
rect 34164 21644 34520 21672
rect 26878 21604 26884 21616
rect 25273 21576 25636 21604
rect 26344 21576 26884 21604
rect 25273 21573 25285 21576
rect 25227 21567 25285 21573
rect 26344 21545 26372 21576
rect 26878 21564 26884 21576
rect 26936 21564 26942 21616
rect 26970 21564 26976 21616
rect 27028 21604 27034 21616
rect 27890 21604 27896 21616
rect 27028 21576 27896 21604
rect 27028 21564 27034 21576
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 28626 21604 28632 21616
rect 28276 21576 28632 21604
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23164 21508 23397 21536
rect 23164 21496 23170 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21505 23719 21539
rect 23661 21499 23719 21505
rect 24581 21539 24639 21545
rect 24581 21505 24593 21539
rect 24627 21536 24639 21539
rect 26329 21539 26387 21545
rect 24627 21508 26280 21536
rect 24627 21505 24639 21508
rect 24581 21499 24639 21505
rect 19116 21440 19472 21468
rect 20901 21471 20959 21477
rect 19116 21428 19122 21440
rect 20901 21437 20913 21471
rect 20947 21468 20959 21471
rect 21174 21468 21180 21480
rect 20947 21440 21180 21468
rect 20947 21437 20959 21440
rect 20901 21431 20959 21437
rect 21174 21428 21180 21440
rect 21232 21468 21238 21480
rect 22646 21468 22652 21480
rect 21232 21440 22652 21468
rect 21232 21428 21238 21440
rect 22646 21428 22652 21440
rect 22704 21428 22710 21480
rect 23676 21468 23704 21499
rect 25774 21468 25780 21480
rect 23676 21440 25780 21468
rect 25774 21428 25780 21440
rect 25832 21428 25838 21480
rect 25866 21428 25872 21480
rect 25924 21468 25930 21480
rect 26145 21471 26203 21477
rect 26145 21468 26157 21471
rect 25924 21440 26157 21468
rect 25924 21428 25930 21440
rect 26145 21437 26157 21440
rect 26191 21437 26203 21471
rect 26252 21468 26280 21508
rect 26329 21505 26341 21539
rect 26375 21505 26387 21539
rect 26329 21499 26387 21505
rect 26421 21539 26479 21545
rect 26421 21505 26433 21539
rect 26467 21536 26479 21539
rect 26467 21508 26648 21536
rect 26467 21505 26479 21508
rect 26421 21499 26479 21505
rect 26510 21468 26516 21480
rect 26252 21440 26516 21468
rect 26145 21431 26203 21437
rect 26510 21428 26516 21440
rect 26568 21428 26574 21480
rect 26620 21468 26648 21508
rect 26694 21496 26700 21548
rect 26752 21536 26758 21548
rect 27157 21539 27215 21545
rect 27157 21536 27169 21539
rect 26752 21508 27169 21536
rect 26752 21496 26758 21508
rect 27157 21505 27169 21508
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21536 27307 21539
rect 28276 21536 28304 21576
rect 28626 21564 28632 21576
rect 28684 21564 28690 21616
rect 30006 21604 30012 21616
rect 29762 21576 30012 21604
rect 30006 21564 30012 21576
rect 30064 21564 30070 21616
rect 30300 21576 31754 21604
rect 30300 21536 30328 21576
rect 30650 21536 30656 21548
rect 27295 21508 28304 21536
rect 29932 21508 30328 21536
rect 30611 21508 30656 21536
rect 27295 21505 27307 21508
rect 27249 21499 27307 21505
rect 29932 21480 29960 21508
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21505 30895 21539
rect 31726 21536 31754 21576
rect 31846 21564 31852 21616
rect 31904 21604 31910 21616
rect 32861 21607 32919 21613
rect 32861 21604 32873 21607
rect 31904 21576 32873 21604
rect 31904 21564 31910 21576
rect 32861 21573 32873 21576
rect 32907 21573 32919 21607
rect 32861 21567 32919 21573
rect 32125 21539 32183 21545
rect 32125 21536 32137 21539
rect 31726 21508 32137 21536
rect 30837 21499 30895 21505
rect 32125 21505 32137 21508
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 32309 21539 32367 21545
rect 32309 21505 32321 21539
rect 32355 21536 32367 21539
rect 32398 21536 32404 21548
rect 32355 21508 32404 21536
rect 32355 21505 32367 21508
rect 32309 21499 32367 21505
rect 28261 21471 28319 21477
rect 26620 21440 27016 21468
rect 10410 21360 10416 21412
rect 10468 21400 10474 21412
rect 10962 21400 10968 21412
rect 10468 21372 10968 21400
rect 10468 21360 10474 21372
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 14550 21360 14556 21412
rect 14608 21360 14614 21412
rect 16117 21403 16175 21409
rect 16117 21369 16129 21403
rect 16163 21400 16175 21403
rect 16850 21400 16856 21412
rect 16163 21372 16856 21400
rect 16163 21369 16175 21372
rect 16117 21363 16175 21369
rect 16850 21360 16856 21372
rect 16908 21360 16914 21412
rect 19426 21360 19432 21412
rect 19484 21400 19490 21412
rect 19613 21403 19671 21409
rect 19613 21400 19625 21403
rect 19484 21372 19625 21400
rect 19484 21360 19490 21372
rect 19613 21369 19625 21372
rect 19659 21369 19671 21403
rect 19613 21363 19671 21369
rect 23290 21360 23296 21412
rect 23348 21400 23354 21412
rect 25406 21400 25412 21412
rect 23348 21372 25412 21400
rect 23348 21360 23354 21372
rect 25406 21360 25412 21372
rect 25464 21360 25470 21412
rect 26418 21360 26424 21412
rect 26476 21400 26482 21412
rect 26988 21409 27016 21440
rect 28261 21437 28273 21471
rect 28307 21437 28319 21471
rect 28534 21468 28540 21480
rect 28495 21440 28540 21468
rect 28261 21431 28319 21437
rect 26973 21403 27031 21409
rect 26476 21372 26521 21400
rect 26476 21360 26482 21372
rect 26973 21369 26985 21403
rect 27019 21369 27031 21403
rect 26973 21363 27031 21369
rect 13814 21332 13820 21344
rect 8864 21304 13820 21332
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 14737 21335 14795 21341
rect 14737 21332 14749 21335
rect 14516 21304 14749 21332
rect 14516 21292 14522 21304
rect 14737 21301 14749 21304
rect 14783 21301 14795 21335
rect 14737 21295 14795 21301
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 16669 21335 16727 21341
rect 16669 21332 16681 21335
rect 16632 21304 16681 21332
rect 16632 21292 16638 21304
rect 16669 21301 16681 21304
rect 16715 21301 16727 21335
rect 16669 21295 16727 21301
rect 18601 21335 18659 21341
rect 18601 21301 18613 21335
rect 18647 21332 18659 21335
rect 18690 21332 18696 21344
rect 18647 21304 18696 21332
rect 18647 21301 18659 21304
rect 18601 21295 18659 21301
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 20349 21335 20407 21341
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20530 21332 20536 21344
rect 20395 21304 20536 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 21082 21292 21088 21344
rect 21140 21332 21146 21344
rect 21269 21335 21327 21341
rect 21269 21332 21281 21335
rect 21140 21304 21281 21332
rect 21140 21292 21146 21304
rect 21269 21301 21281 21304
rect 21315 21301 21327 21335
rect 21269 21295 21327 21301
rect 23385 21335 23443 21341
rect 23385 21301 23397 21335
rect 23431 21332 23443 21335
rect 23750 21332 23756 21344
rect 23431 21304 23756 21332
rect 23431 21301 23443 21304
rect 23385 21295 23443 21301
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 24486 21332 24492 21344
rect 24447 21304 24492 21332
rect 24486 21292 24492 21304
rect 24544 21292 24550 21344
rect 26142 21292 26148 21344
rect 26200 21332 26206 21344
rect 28276 21332 28304 21431
rect 28534 21428 28540 21440
rect 28592 21428 28598 21480
rect 28626 21428 28632 21480
rect 28684 21468 28690 21480
rect 29914 21468 29920 21480
rect 28684 21440 29920 21468
rect 28684 21428 28690 21440
rect 29914 21428 29920 21440
rect 29972 21428 29978 21480
rect 30852 21468 30880 21499
rect 32398 21496 32404 21508
rect 32456 21496 32462 21548
rect 32953 21539 33011 21545
rect 32953 21505 32965 21539
rect 32999 21505 33011 21539
rect 33226 21536 33232 21548
rect 33187 21508 33232 21536
rect 32953 21499 33011 21505
rect 30024 21440 30880 21468
rect 26200 21304 28304 21332
rect 26200 21292 26206 21304
rect 29730 21292 29736 21344
rect 29788 21332 29794 21344
rect 30024 21341 30052 21440
rect 30469 21403 30527 21409
rect 30469 21369 30481 21403
rect 30515 21400 30527 21403
rect 31110 21400 31116 21412
rect 30515 21372 31116 21400
rect 30515 21369 30527 21372
rect 30469 21363 30527 21369
rect 31110 21360 31116 21372
rect 31168 21360 31174 21412
rect 32968 21400 32996 21499
rect 33226 21496 33232 21508
rect 33284 21496 33290 21548
rect 33410 21536 33416 21548
rect 33371 21508 33416 21536
rect 33410 21496 33416 21508
rect 33468 21496 33474 21548
rect 33689 21539 33747 21545
rect 33689 21505 33701 21539
rect 33735 21536 33747 21539
rect 34054 21536 34060 21548
rect 33735 21508 34060 21536
rect 33735 21505 33747 21508
rect 33689 21499 33747 21505
rect 34054 21496 34060 21508
rect 34112 21496 34118 21548
rect 34164 21545 34192 21644
rect 34514 21632 34520 21644
rect 34572 21672 34578 21684
rect 35802 21672 35808 21684
rect 34572 21644 35808 21672
rect 34572 21632 34578 21644
rect 35802 21632 35808 21644
rect 35860 21632 35866 21684
rect 34698 21564 34704 21616
rect 34756 21604 34762 21616
rect 35069 21607 35127 21613
rect 35069 21604 35081 21607
rect 34756 21576 35081 21604
rect 34756 21564 34762 21576
rect 35069 21573 35081 21576
rect 35115 21573 35127 21607
rect 35069 21567 35127 21573
rect 36078 21564 36084 21616
rect 36136 21564 36142 21616
rect 34149 21539 34207 21545
rect 34149 21505 34161 21539
rect 34195 21505 34207 21539
rect 34149 21499 34207 21505
rect 37550 21496 37556 21548
rect 37608 21536 37614 21548
rect 37645 21539 37703 21545
rect 37645 21536 37657 21539
rect 37608 21508 37657 21536
rect 37608 21496 37614 21508
rect 37645 21505 37657 21508
rect 37691 21505 37703 21539
rect 37645 21499 37703 21505
rect 33042 21428 33048 21480
rect 33100 21468 33106 21480
rect 34793 21471 34851 21477
rect 34793 21468 34805 21471
rect 33100 21440 34805 21468
rect 33100 21428 33106 21440
rect 34793 21437 34805 21440
rect 34839 21437 34851 21471
rect 34793 21431 34851 21437
rect 34514 21400 34520 21412
rect 32968 21372 34520 21400
rect 34514 21360 34520 21372
rect 34572 21360 34578 21412
rect 30009 21335 30067 21341
rect 30009 21332 30021 21335
rect 29788 21304 30021 21332
rect 29788 21292 29794 21304
rect 30009 21301 30021 21304
rect 30055 21301 30067 21335
rect 31018 21332 31024 21344
rect 30979 21304 31024 21332
rect 30009 21295 30067 21301
rect 31018 21292 31024 21304
rect 31076 21292 31082 21344
rect 32214 21332 32220 21344
rect 32175 21304 32220 21332
rect 32214 21292 32220 21304
rect 32272 21292 32278 21344
rect 34241 21335 34299 21341
rect 34241 21301 34253 21335
rect 34287 21332 34299 21335
rect 34606 21332 34612 21344
rect 34287 21304 34612 21332
rect 34287 21301 34299 21304
rect 34241 21295 34299 21301
rect 34606 21292 34612 21304
rect 34664 21292 34670 21344
rect 36541 21335 36599 21341
rect 36541 21301 36553 21335
rect 36587 21332 36599 21335
rect 37274 21332 37280 21344
rect 36587 21304 37280 21332
rect 36587 21301 36599 21304
rect 36541 21295 36599 21301
rect 37274 21292 37280 21304
rect 37332 21292 37338 21344
rect 37737 21335 37795 21341
rect 37737 21301 37749 21335
rect 37783 21332 37795 21335
rect 37918 21332 37924 21344
rect 37783 21304 37924 21332
rect 37783 21301 37795 21304
rect 37737 21295 37795 21301
rect 37918 21292 37924 21304
rect 37976 21292 37982 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 5353 21131 5411 21137
rect 5353 21097 5365 21131
rect 5399 21128 5411 21131
rect 5442 21128 5448 21140
rect 5399 21100 5448 21128
rect 5399 21097 5411 21100
rect 5353 21091 5411 21097
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 6365 21131 6423 21137
rect 6365 21097 6377 21131
rect 6411 21128 6423 21131
rect 6546 21128 6552 21140
rect 6411 21100 6552 21128
rect 6411 21097 6423 21100
rect 6365 21091 6423 21097
rect 6546 21088 6552 21100
rect 6604 21088 6610 21140
rect 8205 21131 8263 21137
rect 8205 21097 8217 21131
rect 8251 21128 8263 21131
rect 8386 21128 8392 21140
rect 8251 21100 8392 21128
rect 8251 21097 8263 21100
rect 8205 21091 8263 21097
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 10502 21128 10508 21140
rect 10463 21100 10508 21128
rect 10502 21088 10508 21100
rect 10560 21088 10566 21140
rect 11146 21128 11152 21140
rect 10612 21100 11152 21128
rect 6638 21060 6644 21072
rect 5092 21032 6644 21060
rect 1394 20884 1400 20936
rect 1452 20924 1458 20936
rect 5092 20933 5120 21032
rect 5902 20992 5908 21004
rect 5863 20964 5908 20992
rect 5902 20952 5908 20964
rect 5960 20952 5966 21004
rect 6196 21001 6224 21032
rect 6638 21020 6644 21032
rect 6696 21020 6702 21072
rect 7834 21020 7840 21072
rect 7892 21060 7898 21072
rect 9401 21063 9459 21069
rect 9401 21060 9413 21063
rect 7892 21032 9413 21060
rect 7892 21020 7898 21032
rect 9401 21029 9413 21032
rect 9447 21029 9459 21063
rect 10612 21060 10640 21100
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 13357 21131 13415 21137
rect 13357 21097 13369 21131
rect 13403 21128 13415 21131
rect 13814 21128 13820 21140
rect 13403 21100 13820 21128
rect 13403 21097 13415 21100
rect 13357 21091 13415 21097
rect 13814 21088 13820 21100
rect 13872 21128 13878 21140
rect 14826 21128 14832 21140
rect 13872 21100 14832 21128
rect 13872 21088 13878 21100
rect 14826 21088 14832 21100
rect 14884 21088 14890 21140
rect 20070 21128 20076 21140
rect 19352 21100 20076 21128
rect 9401 21023 9459 21029
rect 10060 21032 10640 21060
rect 10704 21032 11652 21060
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20961 6239 20995
rect 6656 20992 6684 21020
rect 6656 20964 9260 20992
rect 6181 20955 6239 20961
rect 1581 20927 1639 20933
rect 1581 20924 1593 20927
rect 1452 20896 1593 20924
rect 1452 20884 1458 20896
rect 1581 20893 1593 20896
rect 1627 20893 1639 20927
rect 1581 20887 1639 20893
rect 5077 20927 5135 20933
rect 5077 20893 5089 20927
rect 5123 20893 5135 20927
rect 5077 20887 5135 20893
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20924 5411 20927
rect 5994 20924 6000 20936
rect 5399 20896 6000 20924
rect 5399 20893 5411 20896
rect 5353 20887 5411 20893
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 6089 20927 6147 20933
rect 6089 20893 6101 20927
rect 6135 20924 6147 20927
rect 6454 20924 6460 20936
rect 6135 20896 6460 20924
rect 6135 20893 6147 20896
rect 6089 20887 6147 20893
rect 5261 20859 5319 20865
rect 5261 20825 5273 20859
rect 5307 20856 5319 20859
rect 6104 20856 6132 20887
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 6730 20884 6736 20936
rect 6788 20924 6794 20936
rect 6825 20927 6883 20933
rect 6825 20924 6837 20927
rect 6788 20896 6837 20924
rect 6788 20884 6794 20896
rect 6825 20893 6837 20896
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20893 7159 20927
rect 7101 20887 7159 20893
rect 5307 20828 6132 20856
rect 5307 20825 5319 20828
rect 5261 20819 5319 20825
rect 5994 20748 6000 20800
rect 6052 20788 6058 20800
rect 6730 20788 6736 20800
rect 6052 20760 6736 20788
rect 6052 20748 6058 20760
rect 6730 20748 6736 20760
rect 6788 20788 6794 20800
rect 7116 20788 7144 20887
rect 8110 20884 8116 20936
rect 8168 20924 8174 20936
rect 9232 20933 9260 20964
rect 10060 20933 10088 21032
rect 10704 20992 10732 21032
rect 10612 20964 10732 20992
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8168 20896 8953 20924
rect 8168 20884 8174 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 9217 20927 9275 20933
rect 9217 20893 9229 20927
rect 9263 20893 9275 20927
rect 9217 20887 9275 20893
rect 9861 20927 9919 20933
rect 9861 20893 9873 20927
rect 9907 20893 9919 20927
rect 9861 20887 9919 20893
rect 10045 20927 10103 20933
rect 10045 20893 10057 20927
rect 10091 20893 10103 20927
rect 10612 20926 10640 20964
rect 10778 20952 10784 21004
rect 10836 20992 10842 21004
rect 11146 20992 11152 21004
rect 10836 20964 10916 20992
rect 11107 20964 11152 20992
rect 10836 20952 10842 20964
rect 10888 20933 10916 20964
rect 11146 20952 11152 20964
rect 11204 20992 11210 21004
rect 11624 21001 11652 21032
rect 11609 20995 11667 21001
rect 11204 20964 11376 20992
rect 11204 20952 11210 20964
rect 10689 20927 10747 20933
rect 10689 20926 10701 20927
rect 10612 20898 10701 20926
rect 10045 20887 10103 20893
rect 10689 20893 10701 20898
rect 10735 20893 10747 20927
rect 10689 20887 10747 20893
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20893 10931 20927
rect 10873 20887 10931 20893
rect 8294 20856 8300 20868
rect 8255 20828 8300 20856
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 9033 20791 9091 20797
rect 9033 20788 9045 20791
rect 6788 20760 9045 20788
rect 6788 20748 6794 20760
rect 9033 20757 9045 20760
rect 9079 20757 9091 20791
rect 9876 20788 9904 20887
rect 10962 20884 10968 20936
rect 11020 20933 11026 20936
rect 11020 20927 11049 20933
rect 11037 20893 11049 20927
rect 11348 20924 11376 20964
rect 11609 20961 11621 20995
rect 11655 20961 11667 20995
rect 12805 20995 12863 21001
rect 11609 20955 11667 20961
rect 11900 20964 12664 20992
rect 11793 20927 11851 20933
rect 11793 20924 11805 20927
rect 11348 20896 11805 20924
rect 11020 20887 11049 20893
rect 11793 20893 11805 20896
rect 11839 20893 11851 20927
rect 11793 20887 11851 20893
rect 11020 20884 11026 20887
rect 9953 20859 10011 20865
rect 9953 20825 9965 20859
rect 9999 20856 10011 20859
rect 10781 20859 10839 20865
rect 10781 20856 10793 20859
rect 9999 20828 10793 20856
rect 9999 20825 10011 20828
rect 9953 20819 10011 20825
rect 10781 20825 10793 20828
rect 10827 20856 10839 20859
rect 11330 20856 11336 20868
rect 10827 20828 11336 20856
rect 10827 20825 10839 20828
rect 10781 20819 10839 20825
rect 11330 20816 11336 20828
rect 11388 20856 11394 20868
rect 11900 20856 11928 20964
rect 12636 20933 12664 20964
rect 12805 20961 12817 20995
rect 12851 20992 12863 20995
rect 13998 20992 14004 21004
rect 12851 20964 14004 20992
rect 12851 20961 12863 20964
rect 12805 20955 12863 20961
rect 13998 20952 14004 20964
rect 14056 20952 14062 21004
rect 16390 20952 16396 21004
rect 16448 20992 16454 21004
rect 16761 20995 16819 21001
rect 16761 20992 16773 20995
rect 16448 20964 16773 20992
rect 16448 20952 16454 20964
rect 16761 20961 16773 20964
rect 16807 20961 16819 20995
rect 16761 20955 16819 20961
rect 18230 20952 18236 21004
rect 18288 20992 18294 21004
rect 18509 20995 18567 21001
rect 18509 20992 18521 20995
rect 18288 20964 18521 20992
rect 18288 20952 18294 20964
rect 18509 20961 18521 20964
rect 18555 20961 18567 20995
rect 18509 20955 18567 20961
rect 19352 20936 19380 21100
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 21174 21128 21180 21140
rect 21135 21100 21180 21128
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 25887 21131 25945 21137
rect 25887 21097 25899 21131
rect 25933 21128 25945 21131
rect 26234 21128 26240 21140
rect 25933 21100 26240 21128
rect 25933 21097 25945 21100
rect 25887 21091 25945 21097
rect 26234 21088 26240 21100
rect 26292 21088 26298 21140
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 26605 21131 26663 21137
rect 26605 21128 26617 21131
rect 26384 21100 26617 21128
rect 26384 21088 26390 21100
rect 26605 21097 26617 21100
rect 26651 21097 26663 21131
rect 26605 21091 26663 21097
rect 26712 21100 27844 21128
rect 19426 21020 19432 21072
rect 19484 21020 19490 21072
rect 19444 20992 19472 21020
rect 22925 20995 22983 21001
rect 19444 20964 19656 20992
rect 12621 20927 12679 20933
rect 12621 20893 12633 20927
rect 12667 20893 12679 20927
rect 12621 20887 12679 20893
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20924 14151 20927
rect 14734 20924 14740 20936
rect 14139 20896 14740 20924
rect 14139 20893 14151 20896
rect 14093 20887 14151 20893
rect 14734 20884 14740 20896
rect 14792 20884 14798 20936
rect 16485 20927 16543 20933
rect 16485 20893 16497 20927
rect 16531 20924 16543 20927
rect 16574 20924 16580 20936
rect 16531 20896 16580 20924
rect 16531 20893 16543 20896
rect 16485 20887 16543 20893
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 19334 20924 19340 20936
rect 19247 20896 19340 20924
rect 19334 20884 19340 20896
rect 19392 20924 19398 20936
rect 19628 20933 19656 20964
rect 22925 20961 22937 20995
rect 22971 20992 22983 20995
rect 23566 20992 23572 21004
rect 22971 20964 23572 20992
rect 22971 20961 22983 20964
rect 22925 20955 22983 20961
rect 23566 20952 23572 20964
rect 23624 20952 23630 21004
rect 23661 20995 23719 21001
rect 23661 20961 23673 20995
rect 23707 20992 23719 20995
rect 23842 20992 23848 21004
rect 23707 20964 23848 20992
rect 23707 20961 23719 20964
rect 23661 20955 23719 20961
rect 23842 20952 23848 20964
rect 23900 20992 23906 21004
rect 24578 20992 24584 21004
rect 23900 20964 24584 20992
rect 23900 20952 23906 20964
rect 24578 20952 24584 20964
rect 24636 20952 24642 21004
rect 25498 20952 25504 21004
rect 25556 20992 25562 21004
rect 26712 20992 26740 21100
rect 27157 21063 27215 21069
rect 27157 21029 27169 21063
rect 27203 21060 27215 21063
rect 27706 21060 27712 21072
rect 27203 21032 27712 21060
rect 27203 21029 27215 21032
rect 27157 21023 27215 21029
rect 27706 21020 27712 21032
rect 27764 21020 27770 21072
rect 27816 21060 27844 21100
rect 27890 21088 27896 21140
rect 27948 21128 27954 21140
rect 28166 21128 28172 21140
rect 27948 21100 28172 21128
rect 27948 21088 27954 21100
rect 28166 21088 28172 21100
rect 28224 21088 28230 21140
rect 28353 21131 28411 21137
rect 28353 21097 28365 21131
rect 28399 21128 28411 21131
rect 28534 21128 28540 21140
rect 28399 21100 28540 21128
rect 28399 21097 28411 21100
rect 28353 21091 28411 21097
rect 28534 21088 28540 21100
rect 28592 21088 28598 21140
rect 30006 21128 30012 21140
rect 29967 21100 30012 21128
rect 30006 21088 30012 21100
rect 30064 21088 30070 21140
rect 30285 21131 30343 21137
rect 30285 21097 30297 21131
rect 30331 21128 30343 21131
rect 33410 21128 33416 21140
rect 30331 21100 33416 21128
rect 30331 21097 30343 21100
rect 30285 21091 30343 21097
rect 33410 21088 33416 21100
rect 33468 21088 33474 21140
rect 33686 21128 33692 21140
rect 33647 21100 33692 21128
rect 33686 21088 33692 21100
rect 33744 21088 33750 21140
rect 33778 21088 33784 21140
rect 33836 21128 33842 21140
rect 34057 21131 34115 21137
rect 34057 21128 34069 21131
rect 33836 21100 34069 21128
rect 33836 21088 33842 21100
rect 34057 21097 34069 21100
rect 34103 21097 34115 21131
rect 34057 21091 34115 21097
rect 30929 21063 30987 21069
rect 27816 21032 29960 21060
rect 25556 20964 26740 20992
rect 25556 20952 25562 20964
rect 26878 20952 26884 21004
rect 26936 20992 26942 21004
rect 27249 20995 27307 21001
rect 27249 20992 27261 20995
rect 26936 20964 27261 20992
rect 26936 20952 26942 20964
rect 27249 20961 27261 20964
rect 27295 20961 27307 20995
rect 28902 20992 28908 21004
rect 27249 20955 27307 20961
rect 28552 20964 28908 20992
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19392 20896 19441 20924
rect 19392 20884 19398 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20924 19763 20927
rect 19978 20924 19984 20936
rect 19751 20896 19984 20924
rect 19751 20893 19763 20896
rect 19705 20887 19763 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 20349 20927 20407 20933
rect 20349 20893 20361 20927
rect 20395 20893 20407 20927
rect 20349 20887 20407 20893
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20924 20591 20927
rect 20898 20924 20904 20936
rect 20579 20896 20904 20924
rect 20579 20893 20591 20896
rect 20533 20887 20591 20893
rect 11388 20828 11928 20856
rect 11977 20859 12035 20865
rect 11388 20816 11394 20828
rect 11977 20825 11989 20859
rect 12023 20856 12035 20859
rect 12802 20856 12808 20868
rect 12023 20828 12808 20856
rect 12023 20825 12035 20828
rect 11977 20819 12035 20825
rect 11992 20788 12020 20819
rect 12802 20816 12808 20828
rect 12860 20816 12866 20868
rect 12894 20816 12900 20868
rect 12952 20856 12958 20868
rect 13449 20859 13507 20865
rect 13449 20856 13461 20859
rect 12952 20828 13461 20856
rect 12952 20816 12958 20828
rect 13449 20825 13461 20828
rect 13495 20856 13507 20859
rect 13538 20856 13544 20868
rect 13495 20828 13544 20856
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 13538 20816 13544 20828
rect 13596 20816 13602 20868
rect 14360 20859 14418 20865
rect 14360 20825 14372 20859
rect 14406 20856 14418 20859
rect 14642 20856 14648 20868
rect 14406 20828 14648 20856
rect 14406 20825 14418 20828
rect 14360 20819 14418 20825
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 14918 20816 14924 20868
rect 14976 20856 14982 20868
rect 18417 20859 18475 20865
rect 14976 20828 18000 20856
rect 14976 20816 14982 20828
rect 9876 20760 12020 20788
rect 9033 20751 9091 20757
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 12492 20760 12537 20788
rect 12492 20748 12498 20760
rect 13998 20748 14004 20800
rect 14056 20788 14062 20800
rect 15473 20791 15531 20797
rect 15473 20788 15485 20791
rect 14056 20760 15485 20788
rect 14056 20748 14062 20760
rect 15473 20757 15485 20760
rect 15519 20788 15531 20791
rect 15562 20788 15568 20800
rect 15519 20760 15568 20788
rect 15519 20757 15531 20760
rect 15473 20751 15531 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 17972 20797 18000 20828
rect 18417 20825 18429 20859
rect 18463 20856 18475 20859
rect 19245 20859 19303 20865
rect 19245 20856 19257 20859
rect 18463 20828 19257 20856
rect 18463 20825 18475 20828
rect 18417 20819 18475 20825
rect 19245 20825 19257 20828
rect 19291 20856 19303 20859
rect 20364 20856 20392 20887
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 23198 20884 23204 20936
rect 23256 20924 23262 20936
rect 23382 20924 23388 20936
rect 23256 20896 23388 20924
rect 23256 20884 23262 20896
rect 23382 20884 23388 20896
rect 23440 20884 23446 20936
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20924 23535 20927
rect 23934 20924 23940 20936
rect 23523 20896 23940 20924
rect 23523 20893 23535 20896
rect 23477 20887 23535 20893
rect 23934 20884 23940 20896
rect 23992 20884 23998 20936
rect 26142 20884 26148 20936
rect 26200 20924 26206 20936
rect 28552 20933 28580 20964
rect 28902 20952 28908 20964
rect 28960 20952 28966 21004
rect 26730 20927 26788 20933
rect 26730 20924 26742 20927
rect 26200 20896 26245 20924
rect 26436 20896 26742 20924
rect 26200 20884 26206 20896
rect 19291 20828 20392 20856
rect 19291 20825 19303 20828
rect 19245 20819 19303 20825
rect 20438 20816 20444 20868
rect 20496 20856 20502 20868
rect 22646 20856 22652 20868
rect 20496 20828 21482 20856
rect 22607 20828 22652 20856
rect 20496 20816 20502 20828
rect 22646 20816 22652 20828
rect 22704 20816 22710 20868
rect 23566 20816 23572 20868
rect 23624 20856 23630 20868
rect 23624 20828 24702 20856
rect 23624 20816 23630 20828
rect 25774 20816 25780 20868
rect 25832 20856 25838 20868
rect 26436 20856 26464 20896
rect 26730 20893 26742 20896
rect 26776 20893 26788 20927
rect 27709 20927 27767 20933
rect 27709 20924 27721 20927
rect 26730 20887 26788 20893
rect 26896 20896 27721 20924
rect 26896 20856 26924 20896
rect 27709 20893 27721 20896
rect 27755 20893 27767 20927
rect 27709 20887 27767 20893
rect 28537 20927 28595 20933
rect 28537 20893 28549 20927
rect 28583 20893 28595 20927
rect 28537 20887 28595 20893
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 29641 20927 29699 20933
rect 29641 20924 29653 20927
rect 28629 20887 28687 20893
rect 28920 20896 29653 20924
rect 25832 20828 26464 20856
rect 26528 20828 26924 20856
rect 25832 20816 25838 20828
rect 17957 20791 18015 20797
rect 17957 20757 17969 20791
rect 18003 20757 18015 20791
rect 17957 20751 18015 20757
rect 18138 20748 18144 20800
rect 18196 20788 18202 20800
rect 18325 20791 18383 20797
rect 18325 20788 18337 20791
rect 18196 20760 18337 20788
rect 18196 20748 18202 20760
rect 18325 20757 18337 20760
rect 18371 20757 18383 20791
rect 18325 20751 18383 20757
rect 20165 20791 20223 20797
rect 20165 20757 20177 20791
rect 20211 20788 20223 20791
rect 20254 20788 20260 20800
rect 20211 20760 20260 20788
rect 20211 20757 20223 20760
rect 20165 20751 20223 20757
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 23658 20788 23664 20800
rect 23619 20760 23664 20788
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 24397 20791 24455 20797
rect 24397 20757 24409 20791
rect 24443 20788 24455 20791
rect 26326 20788 26332 20800
rect 24443 20760 26332 20788
rect 24443 20757 24455 20760
rect 24397 20751 24455 20757
rect 26326 20748 26332 20760
rect 26384 20788 26390 20800
rect 26528 20788 26556 20828
rect 27522 20816 27528 20868
rect 27580 20856 27586 20868
rect 27580 20828 28028 20856
rect 27580 20816 27586 20828
rect 26786 20788 26792 20800
rect 26384 20760 26556 20788
rect 26747 20760 26792 20788
rect 26384 20748 26390 20760
rect 26786 20748 26792 20760
rect 26844 20748 26850 20800
rect 28000 20788 28028 20828
rect 28074 20816 28080 20868
rect 28132 20856 28138 20868
rect 28353 20859 28411 20865
rect 28353 20856 28365 20859
rect 28132 20828 28365 20856
rect 28132 20816 28138 20828
rect 28353 20825 28365 20828
rect 28399 20825 28411 20859
rect 28353 20819 28411 20825
rect 28644 20788 28672 20887
rect 28920 20868 28948 20896
rect 29641 20893 29653 20896
rect 29687 20893 29699 20927
rect 29641 20887 29699 20893
rect 29730 20884 29736 20936
rect 29788 20924 29794 20936
rect 29788 20896 29881 20924
rect 29788 20884 29794 20896
rect 28902 20816 28908 20868
rect 28960 20816 28966 20868
rect 29086 20816 29092 20868
rect 29144 20856 29150 20868
rect 29748 20856 29776 20884
rect 29144 20828 29776 20856
rect 29144 20816 29150 20828
rect 28000 20760 28672 20788
rect 29932 20788 29960 21032
rect 30929 21029 30941 21063
rect 30975 21060 30987 21063
rect 31110 21060 31116 21072
rect 30975 21032 31116 21060
rect 30975 21029 30987 21032
rect 30929 21023 30987 21029
rect 31110 21020 31116 21032
rect 31168 21020 31174 21072
rect 35621 21063 35679 21069
rect 35621 21060 35633 21063
rect 34164 21032 35633 21060
rect 32030 20952 32036 21004
rect 32088 20992 32094 21004
rect 32677 20995 32735 21001
rect 32677 20992 32689 20995
rect 32088 20964 32689 20992
rect 32088 20952 32094 20964
rect 32677 20961 32689 20964
rect 32723 20992 32735 20995
rect 33042 20992 33048 21004
rect 32723 20964 33048 20992
rect 32723 20961 32735 20964
rect 32677 20955 32735 20961
rect 33042 20952 33048 20964
rect 33100 20952 33106 21004
rect 34164 21001 34192 21032
rect 35621 21029 35633 21032
rect 35667 21060 35679 21063
rect 35710 21060 35716 21072
rect 35667 21032 35716 21060
rect 35667 21029 35679 21032
rect 35621 21023 35679 21029
rect 35710 21020 35716 21032
rect 35768 21020 35774 21072
rect 34149 20995 34207 21001
rect 34149 20961 34161 20995
rect 34195 20961 34207 20995
rect 36446 20992 36452 21004
rect 36407 20964 36452 20992
rect 34149 20955 34207 20961
rect 36446 20952 36452 20964
rect 36504 20952 36510 21004
rect 38102 20992 38108 21004
rect 38063 20964 38108 20992
rect 38102 20952 38108 20964
rect 38160 20952 38166 21004
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20924 30159 20927
rect 30834 20924 30840 20936
rect 30147 20896 30840 20924
rect 30147 20893 30159 20896
rect 30101 20887 30159 20893
rect 30834 20884 30840 20896
rect 30892 20884 30898 20936
rect 33134 20884 33140 20936
rect 33192 20924 33198 20936
rect 33873 20927 33931 20933
rect 33873 20924 33885 20927
rect 33192 20896 33885 20924
rect 33192 20884 33198 20896
rect 33873 20893 33885 20896
rect 33919 20893 33931 20927
rect 36265 20927 36323 20933
rect 36265 20924 36277 20927
rect 33873 20887 33931 20893
rect 34256 20896 36277 20924
rect 31938 20816 31944 20868
rect 31996 20816 32002 20868
rect 32401 20859 32459 20865
rect 32401 20825 32413 20859
rect 32447 20856 32459 20859
rect 33410 20856 33416 20868
rect 32447 20828 33416 20856
rect 32447 20825 32459 20828
rect 32401 20819 32459 20825
rect 33410 20816 33416 20828
rect 33468 20816 33474 20868
rect 34256 20788 34284 20896
rect 36265 20893 36277 20896
rect 36311 20893 36323 20927
rect 36265 20887 36323 20893
rect 35342 20856 35348 20868
rect 35303 20828 35348 20856
rect 35342 20816 35348 20828
rect 35400 20816 35406 20868
rect 35437 20859 35495 20865
rect 35437 20825 35449 20859
rect 35483 20856 35495 20859
rect 37274 20856 37280 20868
rect 35483 20828 37280 20856
rect 35483 20825 35495 20828
rect 35437 20819 35495 20825
rect 37274 20816 37280 20828
rect 37332 20816 37338 20868
rect 29932 20760 34284 20788
rect 34698 20748 34704 20800
rect 34756 20788 34762 20800
rect 35069 20791 35127 20797
rect 35069 20788 35081 20791
rect 34756 20760 35081 20788
rect 34756 20748 34762 20760
rect 35069 20757 35081 20760
rect 35115 20757 35127 20791
rect 35069 20751 35127 20757
rect 35253 20791 35311 20797
rect 35253 20757 35265 20791
rect 35299 20788 35311 20791
rect 35894 20788 35900 20800
rect 35299 20760 35900 20788
rect 35299 20757 35311 20760
rect 35253 20751 35311 20757
rect 35894 20748 35900 20760
rect 35952 20788 35958 20800
rect 36722 20788 36728 20800
rect 35952 20760 36728 20788
rect 35952 20748 35958 20760
rect 36722 20748 36728 20760
rect 36780 20748 36786 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 5813 20587 5871 20593
rect 5813 20553 5825 20587
rect 5859 20584 5871 20587
rect 6638 20584 6644 20596
rect 5859 20556 6644 20584
rect 5859 20553 5871 20556
rect 5813 20547 5871 20553
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 9033 20587 9091 20593
rect 9033 20584 9045 20587
rect 6748 20556 9045 20584
rect 6178 20516 6184 20528
rect 2056 20488 6184 20516
rect 2056 20460 2084 20488
rect 6178 20476 6184 20488
rect 6236 20476 6242 20528
rect 6748 20525 6776 20556
rect 9033 20553 9045 20556
rect 9079 20553 9091 20587
rect 9033 20547 9091 20553
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11701 20587 11759 20593
rect 11701 20584 11713 20587
rect 11572 20556 11713 20584
rect 11572 20544 11578 20556
rect 11701 20553 11713 20556
rect 11747 20553 11759 20587
rect 13630 20584 13636 20596
rect 13591 20556 13636 20584
rect 11701 20547 11759 20553
rect 13630 20544 13636 20556
rect 13688 20544 13694 20596
rect 14642 20544 14648 20596
rect 14700 20584 14706 20596
rect 14737 20587 14795 20593
rect 14737 20584 14749 20587
rect 14700 20556 14749 20584
rect 14700 20544 14706 20556
rect 14737 20553 14749 20556
rect 14783 20553 14795 20587
rect 14737 20547 14795 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16869 20587 16927 20593
rect 16869 20584 16881 20587
rect 15896 20556 16881 20584
rect 15896 20544 15902 20556
rect 16869 20553 16881 20556
rect 16915 20553 16927 20587
rect 16869 20547 16927 20553
rect 18322 20544 18328 20596
rect 18380 20584 18386 20596
rect 19978 20584 19984 20596
rect 18380 20556 19984 20584
rect 18380 20544 18386 20556
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 21821 20587 21879 20593
rect 21821 20553 21833 20587
rect 21867 20584 21879 20587
rect 22646 20584 22652 20596
rect 21867 20556 22652 20584
rect 21867 20553 21879 20556
rect 21821 20547 21879 20553
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 22833 20587 22891 20593
rect 22833 20553 22845 20587
rect 22879 20584 22891 20587
rect 26421 20587 26479 20593
rect 22879 20556 23796 20584
rect 22879 20553 22891 20556
rect 22833 20547 22891 20553
rect 6733 20519 6791 20525
rect 6733 20485 6745 20519
rect 6779 20485 6791 20519
rect 6733 20479 6791 20485
rect 6822 20476 6828 20528
rect 6880 20525 6886 20528
rect 6880 20519 6909 20525
rect 6897 20485 6909 20519
rect 6880 20479 6909 20485
rect 6880 20476 6886 20479
rect 7098 20476 7104 20528
rect 7156 20516 7162 20528
rect 8665 20519 8723 20525
rect 8665 20516 8677 20519
rect 7156 20488 8677 20516
rect 7156 20476 7162 20488
rect 8665 20485 8677 20488
rect 8711 20485 8723 20519
rect 8665 20479 8723 20485
rect 8754 20476 8760 20528
rect 8812 20516 8818 20528
rect 8849 20519 8907 20525
rect 8849 20516 8861 20519
rect 8812 20488 8861 20516
rect 8812 20476 8818 20488
rect 8849 20485 8861 20488
rect 8895 20485 8907 20519
rect 9490 20516 9496 20528
rect 9451 20488 9496 20516
rect 8849 20479 8907 20485
rect 9490 20476 9496 20488
rect 9548 20516 9554 20528
rect 10962 20516 10968 20528
rect 9548 20488 10968 20516
rect 9548 20476 9554 20488
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 11146 20476 11152 20528
rect 11204 20516 11210 20528
rect 12894 20516 12900 20528
rect 11204 20488 12900 20516
rect 11204 20476 11210 20488
rect 12894 20476 12900 20488
rect 12952 20476 12958 20528
rect 13354 20476 13360 20528
rect 13412 20516 13418 20528
rect 14231 20519 14289 20525
rect 14231 20516 14243 20519
rect 13412 20488 14243 20516
rect 13412 20476 13418 20488
rect 14231 20485 14243 20488
rect 14277 20485 14289 20519
rect 14458 20516 14464 20528
rect 14419 20488 14464 20516
rect 14231 20479 14289 20485
rect 14458 20476 14464 20488
rect 14516 20476 14522 20528
rect 15102 20476 15108 20528
rect 15160 20516 15166 20528
rect 15349 20519 15407 20525
rect 15349 20516 15361 20519
rect 15160 20488 15361 20516
rect 15160 20476 15166 20488
rect 15349 20485 15361 20488
rect 15395 20485 15407 20519
rect 15562 20516 15568 20528
rect 15523 20488 15568 20516
rect 15349 20479 15407 20485
rect 15562 20476 15568 20488
rect 15620 20476 15626 20528
rect 16574 20476 16580 20528
rect 16632 20516 16638 20528
rect 16669 20519 16727 20525
rect 16669 20516 16681 20519
rect 16632 20488 16681 20516
rect 16632 20476 16638 20488
rect 16669 20485 16681 20488
rect 16715 20485 16727 20519
rect 18046 20516 18052 20528
rect 17959 20488 18052 20516
rect 16669 20479 16727 20485
rect 2038 20448 2044 20460
rect 1951 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4522 20448 4528 20460
rect 4479 20420 4528 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 4700 20451 4758 20457
rect 4700 20417 4712 20451
rect 4746 20448 4758 20451
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 4746 20420 6377 20448
rect 4746 20417 4758 20420
rect 4700 20411 4758 20417
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6564 20312 6592 20411
rect 6638 20408 6644 20460
rect 6696 20448 6702 20460
rect 7834 20448 7840 20460
rect 6696 20420 6741 20448
rect 7795 20420 7840 20448
rect 6696 20408 6702 20420
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20448 7987 20451
rect 8294 20448 8300 20460
rect 7975 20420 8300 20448
rect 7975 20417 7987 20420
rect 7929 20411 7987 20417
rect 8294 20408 8300 20420
rect 8352 20448 8358 20460
rect 8352 20420 8800 20448
rect 8352 20408 8358 20420
rect 6730 20340 6736 20392
rect 6788 20380 6794 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 6788 20352 7021 20380
rect 6788 20340 6794 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 8110 20380 8116 20392
rect 8071 20352 8116 20380
rect 7009 20343 7067 20349
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 8772 20380 8800 20420
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 9677 20451 9735 20457
rect 9677 20448 9689 20451
rect 9640 20420 9689 20448
rect 9640 20408 9646 20420
rect 9677 20417 9689 20420
rect 9723 20417 9735 20451
rect 10226 20448 10232 20460
rect 10187 20420 10232 20448
rect 9677 20411 9735 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10413 20451 10471 20457
rect 10413 20417 10425 20451
rect 10459 20448 10471 20451
rect 11974 20448 11980 20460
rect 10459 20420 11008 20448
rect 11935 20420 11980 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 9600 20380 9628 20408
rect 10980 20392 11008 20420
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 8772 20352 9628 20380
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 11238 20340 11244 20392
rect 11296 20380 11302 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 11296 20352 11713 20380
rect 11296 20340 11302 20352
rect 11701 20349 11713 20352
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 11885 20383 11943 20389
rect 11885 20349 11897 20383
rect 11931 20380 11943 20383
rect 12434 20380 12440 20392
rect 11931 20352 12440 20380
rect 11931 20349 11943 20352
rect 11885 20343 11943 20349
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 10778 20312 10784 20324
rect 6564 20284 10784 20312
rect 10778 20272 10784 20284
rect 10836 20312 10842 20324
rect 12713 20315 12771 20321
rect 12713 20312 12725 20315
rect 10836 20284 12725 20312
rect 10836 20272 10842 20284
rect 12713 20281 12725 20284
rect 12759 20281 12771 20315
rect 13464 20312 13492 20411
rect 13998 20408 14004 20460
rect 14056 20448 14062 20460
rect 14093 20451 14151 20457
rect 14093 20448 14105 20451
rect 14056 20420 14105 20448
rect 14056 20408 14062 20420
rect 14093 20417 14105 20420
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 14553 20451 14611 20457
rect 14553 20417 14565 20451
rect 14599 20448 14611 20451
rect 15194 20448 15200 20460
rect 14599 20420 15200 20448
rect 14599 20417 14611 20420
rect 14553 20411 14611 20417
rect 14384 20380 14412 20411
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 17972 20457 18000 20488
rect 18046 20476 18052 20488
rect 18104 20516 18110 20528
rect 19426 20516 19432 20528
rect 18104 20488 19432 20516
rect 18104 20476 18110 20488
rect 19426 20476 19432 20488
rect 19484 20476 19490 20528
rect 23658 20516 23664 20528
rect 22296 20488 23664 20516
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20417 18015 20451
rect 18213 20451 18271 20457
rect 18213 20448 18225 20451
rect 17957 20411 18015 20417
rect 18064 20420 18225 20448
rect 14826 20380 14832 20392
rect 14384 20352 14832 20380
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 18064 20380 18092 20420
rect 18213 20417 18225 20420
rect 18259 20417 18271 20451
rect 18213 20411 18271 20417
rect 19150 20408 19156 20460
rect 19208 20448 19214 20460
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 19208 20420 20177 20448
rect 19208 20408 19214 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 19978 20380 19984 20392
rect 17920 20352 18092 20380
rect 19939 20352 19984 20380
rect 17920 20340 17926 20352
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 20070 20340 20076 20392
rect 20128 20380 20134 20392
rect 20128 20352 20173 20380
rect 20128 20340 20134 20352
rect 20254 20340 20260 20392
rect 20312 20380 20318 20392
rect 21284 20380 21312 20411
rect 21818 20408 21824 20460
rect 21876 20448 21882 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21876 20420 22017 20448
rect 21876 20408 21882 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22186 20448 22192 20460
rect 22147 20420 22192 20448
rect 22005 20411 22063 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 22296 20457 22324 20488
rect 23658 20476 23664 20488
rect 23716 20476 23722 20528
rect 23768 20516 23796 20556
rect 26421 20553 26433 20587
rect 26467 20584 26479 20587
rect 26786 20584 26792 20596
rect 26467 20556 26792 20584
rect 26467 20553 26479 20556
rect 26421 20547 26479 20553
rect 26786 20544 26792 20556
rect 26844 20544 26850 20596
rect 27798 20544 27804 20596
rect 27856 20584 27862 20596
rect 27856 20556 27901 20584
rect 27856 20544 27862 20556
rect 28166 20544 28172 20596
rect 28224 20584 28230 20596
rect 28813 20587 28871 20593
rect 28813 20584 28825 20587
rect 28224 20556 28825 20584
rect 28224 20544 28230 20556
rect 28813 20553 28825 20556
rect 28859 20553 28871 20587
rect 33410 20584 33416 20596
rect 33371 20556 33416 20584
rect 28813 20547 28871 20553
rect 33410 20544 33416 20556
rect 33468 20544 33474 20596
rect 34532 20556 37596 20584
rect 23768 20488 24150 20516
rect 28258 20476 28264 20528
rect 28316 20516 28322 20528
rect 28994 20516 29000 20528
rect 28316 20488 29000 20516
rect 28316 20476 28322 20488
rect 28994 20476 29000 20488
rect 29052 20516 29058 20528
rect 29089 20519 29147 20525
rect 29089 20516 29101 20519
rect 29052 20488 29101 20516
rect 29052 20476 29058 20488
rect 29089 20485 29101 20488
rect 29135 20516 29147 20519
rect 30006 20516 30012 20528
rect 29135 20488 30012 20516
rect 29135 20485 29147 20488
rect 29089 20479 29147 20485
rect 30006 20476 30012 20488
rect 30064 20476 30070 20528
rect 32582 20516 32588 20528
rect 30116 20488 32588 20516
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 22741 20451 22799 20457
rect 22741 20448 22753 20451
rect 22704 20420 22753 20448
rect 22704 20408 22710 20420
rect 22741 20417 22753 20420
rect 22787 20448 22799 20451
rect 23290 20448 23296 20460
rect 22787 20420 23296 20448
rect 22787 20417 22799 20420
rect 22741 20411 22799 20417
rect 23290 20408 23296 20420
rect 23348 20408 23354 20460
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26099 20420 27108 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 23382 20380 23388 20392
rect 20312 20352 20357 20380
rect 21284 20352 22094 20380
rect 23343 20352 23388 20380
rect 20312 20340 20318 20352
rect 14918 20312 14924 20324
rect 13464 20284 14924 20312
rect 12713 20275 12771 20281
rect 14918 20272 14924 20284
rect 14976 20272 14982 20324
rect 15102 20272 15108 20324
rect 15160 20312 15166 20324
rect 15197 20315 15255 20321
rect 15197 20312 15209 20315
rect 15160 20284 15209 20312
rect 15160 20272 15166 20284
rect 15197 20281 15209 20284
rect 15243 20281 15255 20315
rect 22066 20312 22094 20352
rect 23382 20340 23388 20352
rect 23440 20340 23446 20392
rect 23661 20383 23719 20389
rect 23661 20349 23673 20383
rect 23707 20380 23719 20383
rect 23750 20380 23756 20392
rect 23707 20352 23756 20380
rect 23707 20349 23719 20352
rect 23661 20343 23719 20349
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 25961 20383 26019 20389
rect 25961 20349 25973 20383
rect 26007 20349 26019 20383
rect 25961 20343 26019 20349
rect 26145 20383 26203 20389
rect 26145 20349 26157 20383
rect 26191 20349 26203 20383
rect 26145 20343 26203 20349
rect 26237 20383 26295 20389
rect 26237 20349 26249 20383
rect 26283 20380 26295 20383
rect 26510 20380 26516 20392
rect 26283 20352 26516 20380
rect 26283 20349 26295 20352
rect 26237 20343 26295 20349
rect 22738 20312 22744 20324
rect 22066 20284 22744 20312
rect 15197 20275 15255 20281
rect 22738 20272 22744 20284
rect 22796 20272 22802 20324
rect 25130 20312 25136 20324
rect 25091 20284 25136 20312
rect 25130 20272 25136 20284
rect 25188 20272 25194 20324
rect 1578 20204 1584 20256
rect 1636 20244 1642 20256
rect 1949 20247 2007 20253
rect 1949 20244 1961 20247
rect 1636 20216 1961 20244
rect 1636 20204 1642 20216
rect 1949 20213 1961 20216
rect 1995 20213 2007 20247
rect 7466 20244 7472 20256
rect 7427 20216 7472 20244
rect 1949 20207 2007 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10413 20247 10471 20253
rect 10413 20244 10425 20247
rect 9824 20216 10425 20244
rect 9824 20204 9830 20216
rect 10413 20213 10425 20216
rect 10459 20213 10471 20247
rect 15378 20244 15384 20256
rect 15339 20216 15384 20244
rect 10413 20207 10471 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 16853 20247 16911 20253
rect 16853 20244 16865 20247
rect 16816 20216 16865 20244
rect 16816 20204 16822 20216
rect 16853 20213 16865 20216
rect 16899 20213 16911 20247
rect 17034 20244 17040 20256
rect 16995 20216 17040 20244
rect 16853 20207 16911 20213
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 19337 20247 19395 20253
rect 19337 20244 19349 20247
rect 18288 20216 19349 20244
rect 18288 20204 18294 20216
rect 19337 20213 19349 20216
rect 19383 20213 19395 20247
rect 19337 20207 19395 20213
rect 19797 20247 19855 20253
rect 19797 20213 19809 20247
rect 19843 20244 19855 20247
rect 19978 20244 19984 20256
rect 19843 20216 19984 20244
rect 19843 20213 19855 20216
rect 19797 20207 19855 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 20806 20204 20812 20256
rect 20864 20244 20870 20256
rect 21085 20247 21143 20253
rect 21085 20244 21097 20247
rect 20864 20216 21097 20244
rect 20864 20204 20870 20216
rect 21085 20213 21097 20216
rect 21131 20244 21143 20247
rect 23842 20244 23848 20256
rect 21131 20216 23848 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 25682 20204 25688 20256
rect 25740 20244 25746 20256
rect 25976 20244 26004 20343
rect 26160 20312 26188 20343
rect 26510 20340 26516 20352
rect 26568 20340 26574 20392
rect 27080 20380 27108 20420
rect 27430 20408 27436 20460
rect 27488 20448 27494 20460
rect 27605 20451 27663 20457
rect 27605 20448 27617 20451
rect 27488 20420 27617 20448
rect 27488 20408 27494 20420
rect 27605 20417 27617 20420
rect 27651 20417 27663 20451
rect 27605 20411 27663 20417
rect 27890 20408 27896 20460
rect 27948 20448 27954 20460
rect 27985 20451 28043 20457
rect 27985 20448 27997 20451
rect 27948 20420 27997 20448
rect 27948 20408 27954 20420
rect 27985 20417 27997 20420
rect 28031 20448 28043 20451
rect 28721 20451 28779 20457
rect 28721 20448 28733 20451
rect 28031 20420 28733 20448
rect 28031 20417 28043 20420
rect 27985 20411 28043 20417
rect 28721 20417 28733 20420
rect 28767 20417 28779 20451
rect 28721 20411 28779 20417
rect 28902 20408 28908 20460
rect 28960 20448 28966 20460
rect 28960 20420 29053 20448
rect 28960 20408 28966 20420
rect 27706 20380 27712 20392
rect 27080 20352 27712 20380
rect 27706 20340 27712 20352
rect 27764 20340 27770 20392
rect 27798 20340 27804 20392
rect 27856 20380 27862 20392
rect 28077 20383 28135 20389
rect 28077 20380 28089 20383
rect 27856 20352 28089 20380
rect 27856 20340 27862 20352
rect 28077 20349 28089 20352
rect 28123 20349 28135 20383
rect 28077 20343 28135 20349
rect 28350 20340 28356 20392
rect 28408 20380 28414 20392
rect 28537 20383 28595 20389
rect 28537 20380 28549 20383
rect 28408 20352 28549 20380
rect 28408 20340 28414 20352
rect 28537 20349 28549 20352
rect 28583 20349 28595 20383
rect 28537 20343 28595 20349
rect 26970 20312 26976 20324
rect 26160 20284 26976 20312
rect 26970 20272 26976 20284
rect 27028 20272 27034 20324
rect 27724 20312 27752 20340
rect 28920 20312 28948 20408
rect 28994 20340 29000 20392
rect 29052 20380 29058 20392
rect 30116 20380 30144 20488
rect 32582 20476 32588 20488
rect 32640 20476 32646 20528
rect 33962 20476 33968 20528
rect 34020 20516 34026 20528
rect 34532 20516 34560 20556
rect 34020 20488 34560 20516
rect 34020 20476 34026 20488
rect 30834 20448 30840 20460
rect 30795 20420 30840 20448
rect 30834 20408 30840 20420
rect 30892 20408 30898 20460
rect 31478 20448 31484 20460
rect 31439 20420 31484 20448
rect 31478 20408 31484 20420
rect 31536 20408 31542 20460
rect 31662 20408 31668 20460
rect 31720 20448 31726 20460
rect 33597 20451 33655 20457
rect 33597 20448 33609 20451
rect 31720 20420 33609 20448
rect 31720 20408 31726 20420
rect 33597 20417 33609 20420
rect 33643 20417 33655 20451
rect 33597 20411 33655 20417
rect 33689 20451 33747 20457
rect 33689 20417 33701 20451
rect 33735 20448 33747 20451
rect 33870 20448 33876 20460
rect 33735 20420 33876 20448
rect 33735 20417 33747 20420
rect 33689 20411 33747 20417
rect 33870 20408 33876 20420
rect 33928 20408 33934 20460
rect 34330 20448 34336 20460
rect 34291 20420 34336 20448
rect 34330 20408 34336 20420
rect 34388 20408 34394 20460
rect 34532 20457 34560 20488
rect 34606 20476 34612 20528
rect 34664 20516 34670 20528
rect 34664 20488 35282 20516
rect 34664 20476 34670 20488
rect 36538 20476 36544 20528
rect 36596 20516 36602 20528
rect 37274 20516 37280 20528
rect 36596 20488 36768 20516
rect 37235 20488 37280 20516
rect 36596 20476 36602 20488
rect 36740 20457 36768 20488
rect 37274 20476 37280 20488
rect 37332 20476 37338 20528
rect 34517 20451 34575 20457
rect 34517 20417 34529 20451
rect 34563 20417 34575 20451
rect 34517 20411 34575 20417
rect 36725 20451 36783 20457
rect 36725 20417 36737 20451
rect 36771 20417 36783 20451
rect 37458 20448 37464 20460
rect 37419 20420 37464 20448
rect 36725 20411 36783 20417
rect 37458 20408 37464 20420
rect 37516 20408 37522 20460
rect 37568 20457 37596 20556
rect 37553 20451 37611 20457
rect 37553 20417 37565 20451
rect 37599 20417 37611 20451
rect 37553 20411 37611 20417
rect 29052 20352 30144 20380
rect 30561 20383 30619 20389
rect 29052 20340 29058 20352
rect 30561 20349 30573 20383
rect 30607 20380 30619 20383
rect 30926 20380 30932 20392
rect 30607 20352 30932 20380
rect 30607 20349 30619 20352
rect 30561 20343 30619 20349
rect 27080 20284 27552 20312
rect 27724 20284 28948 20312
rect 27080 20244 27108 20284
rect 27430 20244 27436 20256
rect 25740 20216 27108 20244
rect 27391 20216 27436 20244
rect 25740 20204 25746 20216
rect 27430 20204 27436 20216
rect 27488 20204 27494 20256
rect 27524 20244 27552 20284
rect 29178 20272 29184 20324
rect 29236 20312 29242 20324
rect 29730 20312 29736 20324
rect 29236 20284 29736 20312
rect 29236 20272 29242 20284
rect 29730 20272 29736 20284
rect 29788 20312 29794 20324
rect 30576 20312 30604 20343
rect 30926 20340 30932 20352
rect 30984 20340 30990 20392
rect 32122 20380 32128 20392
rect 32083 20352 32128 20380
rect 32122 20340 32128 20352
rect 32180 20340 32186 20392
rect 33781 20383 33839 20389
rect 33781 20349 33793 20383
rect 33827 20349 33839 20383
rect 33781 20343 33839 20349
rect 31294 20312 31300 20324
rect 29788 20284 30604 20312
rect 31255 20284 31300 20312
rect 29788 20272 29794 20284
rect 31294 20272 31300 20284
rect 31352 20272 31358 20324
rect 31386 20272 31392 20324
rect 31444 20312 31450 20324
rect 33796 20312 33824 20343
rect 35710 20340 35716 20392
rect 35768 20380 35774 20392
rect 36449 20383 36507 20389
rect 36449 20380 36461 20383
rect 35768 20352 36461 20380
rect 35768 20340 35774 20352
rect 36449 20349 36461 20352
rect 36495 20349 36507 20383
rect 36449 20343 36507 20349
rect 31444 20284 33824 20312
rect 34977 20315 35035 20321
rect 31444 20272 31450 20284
rect 34977 20281 34989 20315
rect 35023 20312 35035 20315
rect 35342 20312 35348 20324
rect 35023 20284 35348 20312
rect 35023 20281 35035 20284
rect 34977 20275 35035 20281
rect 28810 20244 28816 20256
rect 27524 20216 28816 20244
rect 28810 20204 28816 20216
rect 28868 20204 28874 20256
rect 30650 20204 30656 20256
rect 30708 20244 30714 20256
rect 30834 20244 30840 20256
rect 30708 20216 30840 20244
rect 30708 20204 30714 20216
rect 30834 20204 30840 20216
rect 30892 20244 30898 20256
rect 32355 20247 32413 20253
rect 32355 20244 32367 20247
rect 30892 20216 32367 20244
rect 30892 20204 30898 20216
rect 32355 20213 32367 20216
rect 32401 20213 32413 20247
rect 34422 20244 34428 20256
rect 34383 20216 34428 20244
rect 32355 20207 32413 20213
rect 34422 20204 34428 20216
rect 34480 20204 34486 20256
rect 34514 20204 34520 20256
rect 34572 20244 34578 20256
rect 34992 20244 35020 20275
rect 35342 20272 35348 20284
rect 35400 20272 35406 20324
rect 37277 20315 37335 20321
rect 37277 20281 37289 20315
rect 37323 20312 37335 20315
rect 37366 20312 37372 20324
rect 37323 20284 37372 20312
rect 37323 20281 37335 20284
rect 37277 20275 37335 20281
rect 37366 20272 37372 20284
rect 37424 20272 37430 20324
rect 34572 20216 35020 20244
rect 34572 20204 34578 20216
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 6549 20043 6607 20049
rect 6549 20009 6561 20043
rect 6595 20040 6607 20043
rect 6638 20040 6644 20052
rect 6595 20012 6644 20040
rect 6595 20009 6607 20012
rect 6549 20003 6607 20009
rect 6638 20000 6644 20012
rect 6696 20000 6702 20052
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12161 20043 12219 20049
rect 12161 20040 12173 20043
rect 12032 20012 12173 20040
rect 12032 20000 12038 20012
rect 12161 20009 12173 20012
rect 12207 20009 12219 20043
rect 12161 20003 12219 20009
rect 13354 20000 13360 20052
rect 13412 20040 13418 20052
rect 14642 20040 14648 20052
rect 13412 20012 14648 20040
rect 13412 20000 13418 20012
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 15194 20040 15200 20052
rect 15155 20012 15200 20040
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15562 20000 15568 20052
rect 15620 20040 15626 20052
rect 16022 20040 16028 20052
rect 15620 20012 16028 20040
rect 15620 20000 15626 20012
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16209 20043 16267 20049
rect 16209 20040 16221 20043
rect 16172 20012 16221 20040
rect 16172 20000 16178 20012
rect 16209 20009 16221 20012
rect 16255 20009 16267 20043
rect 16209 20003 16267 20009
rect 16298 20000 16304 20052
rect 16356 20040 16362 20052
rect 16761 20043 16819 20049
rect 16761 20040 16773 20043
rect 16356 20012 16773 20040
rect 16356 20000 16362 20012
rect 16761 20009 16773 20012
rect 16807 20040 16819 20043
rect 18322 20040 18328 20052
rect 16807 20012 18328 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18506 20040 18512 20052
rect 18467 20012 18512 20040
rect 18506 20000 18512 20012
rect 18564 20000 18570 20052
rect 19429 20043 19487 20049
rect 19429 20009 19441 20043
rect 19475 20040 19487 20043
rect 20346 20040 20352 20052
rect 19475 20012 20352 20040
rect 19475 20009 19487 20012
rect 19429 20003 19487 20009
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 23106 20040 23112 20052
rect 23067 20012 23112 20040
rect 23106 20000 23112 20012
rect 23164 20000 23170 20052
rect 27062 20000 27068 20052
rect 27120 20040 27126 20052
rect 27249 20043 27307 20049
rect 27249 20040 27261 20043
rect 27120 20012 27261 20040
rect 27120 20000 27126 20012
rect 27249 20009 27261 20012
rect 27295 20009 27307 20043
rect 27249 20003 27307 20009
rect 27433 20043 27491 20049
rect 27433 20009 27445 20043
rect 27479 20040 27491 20043
rect 27522 20040 27528 20052
rect 27479 20012 27528 20040
rect 27479 20009 27491 20012
rect 27433 20003 27491 20009
rect 27522 20000 27528 20012
rect 27580 20000 27586 20052
rect 28902 20000 28908 20052
rect 28960 20040 28966 20052
rect 30098 20040 30104 20052
rect 28960 20012 30104 20040
rect 28960 20000 28966 20012
rect 30098 20000 30104 20012
rect 30156 20000 30162 20052
rect 31297 20043 31355 20049
rect 31297 20009 31309 20043
rect 31343 20040 31355 20043
rect 31386 20040 31392 20052
rect 31343 20012 31392 20040
rect 31343 20009 31355 20012
rect 31297 20003 31355 20009
rect 31386 20000 31392 20012
rect 31444 20000 31450 20052
rect 32306 20000 32312 20052
rect 32364 20040 32370 20052
rect 32677 20043 32735 20049
rect 32677 20040 32689 20043
rect 32364 20012 32689 20040
rect 32364 20000 32370 20012
rect 32677 20009 32689 20012
rect 32723 20009 32735 20043
rect 35710 20040 35716 20052
rect 35671 20012 35716 20040
rect 32677 20003 32735 20009
rect 35710 20000 35716 20012
rect 35768 20000 35774 20052
rect 6454 19972 6460 19984
rect 6367 19944 6460 19972
rect 6454 19932 6460 19944
rect 6512 19972 6518 19984
rect 6512 19944 7420 19972
rect 6512 19932 6518 19944
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 1578 19904 1584 19916
rect 1539 19876 1584 19904
rect 1578 19864 1584 19876
rect 1636 19864 1642 19916
rect 1854 19904 1860 19916
rect 1815 19876 1860 19904
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 6472 19845 6500 19932
rect 7098 19904 7104 19916
rect 7059 19876 7104 19904
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7392 19913 7420 19944
rect 7377 19907 7435 19913
rect 7377 19873 7389 19907
rect 7423 19904 7435 19907
rect 8110 19904 8116 19916
rect 7423 19876 8116 19904
rect 7423 19873 7435 19876
rect 7377 19867 7435 19873
rect 8110 19864 8116 19876
rect 8168 19864 8174 19916
rect 11992 19904 12020 20000
rect 15378 19972 15384 19984
rect 13280 19944 15384 19972
rect 10980 19876 12020 19904
rect 6457 19839 6515 19845
rect 6457 19805 6469 19839
rect 6503 19805 6515 19839
rect 6457 19799 6515 19805
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19836 6699 19839
rect 6730 19836 6736 19848
rect 6687 19808 6736 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 8662 19796 8668 19848
rect 8720 19836 8726 19848
rect 8938 19836 8944 19848
rect 8720 19808 8944 19836
rect 8720 19796 8726 19808
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 9582 19796 9588 19848
rect 9640 19836 9646 19848
rect 10980 19845 11008 19876
rect 13078 19864 13084 19916
rect 13136 19904 13142 19916
rect 13280 19904 13308 19944
rect 15378 19932 15384 19944
rect 15436 19932 15442 19984
rect 16666 19972 16672 19984
rect 15948 19944 16672 19972
rect 13136 19876 13308 19904
rect 13136 19864 13142 19876
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 9640 19808 10977 19836
rect 9640 19796 9646 19808
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11054 19796 11060 19848
rect 11112 19836 11118 19848
rect 11241 19839 11299 19845
rect 11241 19836 11253 19839
rect 11112 19808 11253 19836
rect 11112 19796 11118 19808
rect 11241 19805 11253 19808
rect 11287 19805 11299 19839
rect 13170 19836 13176 19848
rect 13131 19808 13176 19836
rect 11241 19799 11299 19805
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 13280 19845 13308 19876
rect 13541 19907 13599 19913
rect 13541 19873 13553 19907
rect 13587 19904 13599 19907
rect 13722 19904 13728 19916
rect 13587 19876 13728 19904
rect 13587 19873 13599 19876
rect 13541 19867 13599 19873
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 14148 19876 14289 19904
rect 14148 19864 14154 19876
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 14277 19867 14335 19873
rect 14550 19864 14556 19916
rect 14608 19904 14614 19916
rect 15948 19913 15976 19944
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 17310 19932 17316 19984
rect 17368 19972 17374 19984
rect 17368 19944 18644 19972
rect 17368 19932 17374 19944
rect 15933 19907 15991 19913
rect 14608 19876 14653 19904
rect 14608 19864 14614 19876
rect 15933 19873 15945 19907
rect 15979 19873 15991 19907
rect 15933 19867 15991 19873
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 16816 19876 17540 19904
rect 16816 19864 16822 19876
rect 17512 19848 17540 19876
rect 18230 19864 18236 19916
rect 18288 19904 18294 19916
rect 18509 19907 18567 19913
rect 18509 19904 18521 19907
rect 18288 19876 18521 19904
rect 18288 19864 18294 19876
rect 18509 19873 18521 19876
rect 18555 19873 18567 19907
rect 18616 19904 18644 19944
rect 19334 19932 19340 19984
rect 19392 19972 19398 19984
rect 19613 19975 19671 19981
rect 19613 19972 19625 19975
rect 19392 19944 19625 19972
rect 19392 19932 19398 19944
rect 19613 19941 19625 19944
rect 19659 19941 19671 19975
rect 19613 19935 19671 19941
rect 23198 19932 23204 19984
rect 23256 19972 23262 19984
rect 23385 19975 23443 19981
rect 23385 19972 23397 19975
rect 23256 19944 23397 19972
rect 23256 19932 23262 19944
rect 23385 19941 23397 19944
rect 23431 19941 23443 19975
rect 32490 19972 32496 19984
rect 23385 19935 23443 19941
rect 28828 19944 32496 19972
rect 20714 19904 20720 19916
rect 18616 19876 19564 19904
rect 20675 19876 20720 19904
rect 18509 19867 18567 19873
rect 13265 19839 13323 19845
rect 13265 19805 13277 19839
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19836 14519 19839
rect 14642 19836 14648 19848
rect 14507 19808 14648 19836
rect 14507 19805 14519 19808
rect 14461 19799 14519 19805
rect 9030 19728 9036 19780
rect 9088 19768 9094 19780
rect 9186 19771 9244 19777
rect 9186 19768 9198 19771
rect 9088 19740 9198 19768
rect 9088 19728 9094 19740
rect 9186 19737 9198 19740
rect 9232 19737 9244 19771
rect 9186 19731 9244 19737
rect 12253 19771 12311 19777
rect 12253 19737 12265 19771
rect 12299 19768 12311 19771
rect 13078 19768 13084 19780
rect 12299 19740 13084 19768
rect 12299 19737 12311 19740
rect 12253 19731 12311 19737
rect 13078 19728 13084 19740
rect 13136 19728 13142 19780
rect 13538 19728 13544 19780
rect 13596 19768 13602 19780
rect 14384 19768 14412 19799
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19836 15807 19839
rect 15838 19836 15844 19848
rect 15795 19808 15844 19836
rect 15795 19805 15807 19808
rect 15749 19799 15807 19805
rect 13596 19740 14412 19768
rect 13596 19728 13602 19740
rect 15194 19728 15200 19780
rect 15252 19768 15258 19780
rect 15304 19768 15332 19799
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19836 16083 19839
rect 16574 19836 16580 19848
rect 16071 19808 16580 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16850 19836 16856 19848
rect 16811 19808 16856 19836
rect 16669 19799 16727 19805
rect 16684 19768 16712 19799
rect 16850 19796 16856 19808
rect 16908 19796 16914 19848
rect 17218 19836 17224 19848
rect 17179 19808 17224 19836
rect 17218 19796 17224 19808
rect 17276 19796 17282 19848
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 18417 19839 18475 19845
rect 17552 19808 17597 19836
rect 17552 19796 17558 19808
rect 18417 19805 18429 19839
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18739 19833 19288 19836
rect 18739 19808 19380 19833
rect 18739 19805 18751 19808
rect 19260 19805 19380 19808
rect 18693 19799 18751 19805
rect 17126 19768 17132 19780
rect 15252 19740 17132 19768
rect 15252 19728 15258 19740
rect 17126 19728 17132 19740
rect 17184 19728 17190 19780
rect 18432 19768 18460 19799
rect 19150 19768 19156 19780
rect 18432 19740 19156 19768
rect 19150 19728 19156 19740
rect 19208 19728 19214 19780
rect 19245 19771 19303 19777
rect 19245 19737 19257 19771
rect 19291 19737 19303 19771
rect 19245 19731 19303 19737
rect 10318 19700 10324 19712
rect 10279 19672 10324 19700
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 10778 19700 10784 19712
rect 10739 19672 10784 19700
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 11146 19700 11152 19712
rect 11107 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 13354 19700 13360 19712
rect 13315 19672 13360 19700
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13446 19660 13452 19712
rect 13504 19700 13510 19712
rect 13504 19672 13549 19700
rect 13504 19660 13510 19672
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14093 19703 14151 19709
rect 14093 19700 14105 19703
rect 13872 19672 14105 19700
rect 13872 19660 13878 19672
rect 14093 19669 14105 19672
rect 14139 19669 14151 19703
rect 14093 19663 14151 19669
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 18233 19703 18291 19709
rect 18233 19700 18245 19703
rect 15160 19672 18245 19700
rect 15160 19660 15166 19672
rect 18233 19669 18245 19672
rect 18279 19669 18291 19703
rect 18233 19663 18291 19669
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 19260 19700 19288 19731
rect 18380 19672 19288 19700
rect 19352 19700 19380 19805
rect 19445 19771 19503 19777
rect 19445 19737 19457 19771
rect 19491 19768 19503 19771
rect 19536 19768 19564 19876
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 28350 19864 28356 19916
rect 28408 19904 28414 19916
rect 28828 19904 28856 19944
rect 32490 19932 32496 19944
rect 32548 19972 32554 19984
rect 33137 19975 33195 19981
rect 33137 19972 33149 19975
rect 32548 19944 33149 19972
rect 32548 19932 32554 19944
rect 33137 19941 33149 19944
rect 33183 19941 33195 19975
rect 33137 19935 33195 19941
rect 37826 19932 37832 19984
rect 37884 19972 37890 19984
rect 37884 19944 38148 19972
rect 37884 19932 37890 19944
rect 28408 19876 28856 19904
rect 28408 19864 28414 19876
rect 22370 19836 22376 19848
rect 22331 19808 22376 19836
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19805 23351 19839
rect 23474 19836 23480 19848
rect 23435 19808 23480 19836
rect 23293 19799 23351 19805
rect 19491 19740 19564 19768
rect 23308 19768 23336 19799
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19836 23627 19839
rect 24486 19836 24492 19848
rect 23615 19808 24492 19836
rect 23615 19805 23627 19808
rect 23569 19799 23627 19805
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19836 24639 19839
rect 24946 19836 24952 19848
rect 24627 19808 24952 19836
rect 24627 19805 24639 19808
rect 24581 19799 24639 19805
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 25130 19796 25136 19848
rect 25188 19836 25194 19848
rect 25593 19839 25651 19845
rect 25593 19836 25605 19839
rect 25188 19808 25605 19836
rect 25188 19796 25194 19808
rect 25593 19805 25605 19808
rect 25639 19805 25651 19839
rect 25593 19799 25651 19805
rect 25869 19839 25927 19845
rect 25869 19805 25881 19839
rect 25915 19836 25927 19839
rect 26510 19836 26516 19848
rect 25915 19808 26516 19836
rect 25915 19805 25927 19808
rect 25869 19799 25927 19805
rect 26510 19796 26516 19808
rect 26568 19796 26574 19848
rect 28442 19796 28448 19848
rect 28500 19836 28506 19848
rect 28828 19845 28856 19876
rect 28902 19864 28908 19916
rect 28960 19904 28966 19916
rect 29638 19904 29644 19916
rect 28960 19876 29644 19904
rect 28960 19864 28966 19876
rect 29638 19864 29644 19876
rect 29696 19864 29702 19916
rect 31110 19904 31116 19916
rect 31071 19876 31116 19904
rect 31110 19864 31116 19876
rect 31168 19864 31174 19916
rect 32048 19876 33272 19904
rect 32048 19848 32076 19876
rect 28629 19839 28687 19845
rect 28629 19836 28641 19839
rect 28500 19808 28641 19836
rect 28500 19796 28506 19808
rect 28629 19805 28641 19808
rect 28675 19805 28687 19839
rect 28629 19799 28687 19805
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19805 28871 19839
rect 28813 19799 28871 19805
rect 28997 19839 29055 19845
rect 28997 19805 29009 19839
rect 29043 19838 29055 19839
rect 29043 19836 29132 19838
rect 29043 19810 29500 19836
rect 29043 19805 29055 19810
rect 29104 19808 29500 19810
rect 28997 19799 29055 19805
rect 24118 19768 24124 19780
rect 23308 19740 24124 19768
rect 19491 19737 19503 19740
rect 19445 19731 19503 19737
rect 24118 19728 24124 19740
rect 24176 19728 24182 19780
rect 27430 19777 27436 19780
rect 27417 19771 27436 19777
rect 27417 19737 27429 19771
rect 27417 19731 27436 19737
rect 27430 19728 27436 19731
rect 27488 19728 27494 19780
rect 27614 19768 27620 19780
rect 27575 19740 27620 19768
rect 27614 19728 27620 19740
rect 27672 19728 27678 19780
rect 29472 19768 29500 19808
rect 29546 19796 29552 19848
rect 29604 19836 29610 19848
rect 29604 19808 29649 19836
rect 29604 19796 29610 19808
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30009 19839 30067 19845
rect 30009 19838 30021 19839
rect 29788 19808 29833 19836
rect 29932 19810 30021 19838
rect 29788 19796 29794 19808
rect 29822 19768 29828 19780
rect 29472 19740 29828 19768
rect 20898 19700 20904 19712
rect 19352 19672 20904 19700
rect 18380 19660 18386 19672
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 23842 19660 23848 19712
rect 23900 19700 23906 19712
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 23900 19672 24409 19700
rect 23900 19660 23906 19672
rect 24397 19669 24409 19672
rect 24443 19669 24455 19703
rect 24397 19663 24455 19669
rect 27706 19660 27712 19712
rect 27764 19700 27770 19712
rect 28966 19711 29224 19739
rect 29822 19728 29828 19740
rect 29880 19768 29886 19780
rect 29932 19768 29960 19810
rect 30009 19805 30021 19810
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 30558 19796 30564 19848
rect 30616 19836 30622 19848
rect 30653 19839 30711 19845
rect 30653 19836 30665 19839
rect 30616 19808 30665 19836
rect 30616 19796 30622 19808
rect 30653 19805 30665 19808
rect 30699 19805 30711 19839
rect 30653 19799 30711 19805
rect 30834 19796 30840 19848
rect 30892 19836 30898 19848
rect 31021 19839 31079 19845
rect 31021 19836 31033 19839
rect 30892 19808 31033 19836
rect 30892 19796 30898 19808
rect 31021 19805 31033 19808
rect 31067 19805 31079 19839
rect 32030 19836 32036 19848
rect 31943 19808 32036 19836
rect 31021 19799 31079 19805
rect 32030 19796 32036 19808
rect 32088 19796 32094 19848
rect 32214 19836 32220 19848
rect 32175 19808 32220 19836
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 32309 19839 32367 19845
rect 32309 19805 32321 19839
rect 32355 19805 32367 19839
rect 32309 19799 32367 19805
rect 32401 19839 32459 19845
rect 32401 19805 32413 19839
rect 32447 19836 32459 19839
rect 32950 19836 32956 19848
rect 32447 19808 32956 19836
rect 32447 19805 32459 19808
rect 32401 19799 32459 19805
rect 29880 19740 29960 19768
rect 29880 19728 29886 19740
rect 31662 19728 31668 19780
rect 31720 19768 31726 19780
rect 32324 19768 32352 19799
rect 32950 19796 32956 19808
rect 33008 19796 33014 19848
rect 31720 19740 32352 19768
rect 33244 19768 33272 19876
rect 34422 19864 34428 19916
rect 34480 19904 34486 19916
rect 37090 19904 37096 19916
rect 34480 19876 35296 19904
rect 37051 19876 37096 19904
rect 34480 19864 34486 19876
rect 33410 19836 33416 19848
rect 33323 19808 33416 19836
rect 33410 19796 33416 19808
rect 33468 19836 33474 19848
rect 34698 19836 34704 19848
rect 33468 19808 34704 19836
rect 33468 19796 33474 19808
rect 34698 19796 34704 19808
rect 34756 19796 34762 19848
rect 34974 19796 34980 19848
rect 35032 19836 35038 19848
rect 35268 19845 35296 19876
rect 37090 19864 37096 19876
rect 37148 19864 37154 19916
rect 37918 19904 37924 19916
rect 37879 19876 37924 19904
rect 37918 19864 37924 19876
rect 37976 19864 37982 19916
rect 38120 19913 38148 19944
rect 38105 19907 38163 19913
rect 38105 19873 38117 19907
rect 38151 19873 38163 19907
rect 38105 19867 38163 19873
rect 35069 19839 35127 19845
rect 35069 19836 35081 19839
rect 35032 19808 35081 19836
rect 35032 19796 35038 19808
rect 35069 19805 35081 19808
rect 35115 19805 35127 19839
rect 35069 19799 35127 19805
rect 35253 19839 35311 19845
rect 35253 19805 35265 19839
rect 35299 19805 35311 19839
rect 35253 19799 35311 19805
rect 35345 19839 35403 19845
rect 35345 19805 35357 19839
rect 35391 19805 35403 19839
rect 35345 19799 35403 19805
rect 34992 19768 35020 19796
rect 33244 19740 35020 19768
rect 35360 19768 35388 19799
rect 35434 19796 35440 19848
rect 35492 19836 35498 19848
rect 35492 19808 35537 19836
rect 35492 19796 35498 19808
rect 35526 19768 35532 19780
rect 35360 19740 35532 19768
rect 31720 19728 31726 19740
rect 35526 19728 35532 19740
rect 35584 19728 35590 19780
rect 28966 19700 28994 19711
rect 27764 19672 28994 19700
rect 29196 19700 29224 19711
rect 29917 19703 29975 19709
rect 29917 19700 29929 19703
rect 29196 19672 29929 19700
rect 27764 19660 27770 19672
rect 29917 19669 29929 19672
rect 29963 19669 29975 19703
rect 29917 19663 29975 19669
rect 30650 19660 30656 19712
rect 30708 19700 30714 19712
rect 30745 19703 30803 19709
rect 30745 19700 30757 19703
rect 30708 19672 30757 19700
rect 30708 19660 30714 19672
rect 30745 19669 30757 19672
rect 30791 19669 30803 19703
rect 30926 19700 30932 19712
rect 30887 19672 30932 19700
rect 30745 19663 30803 19669
rect 30926 19660 30932 19672
rect 30984 19660 30990 19712
rect 33318 19700 33324 19712
rect 33279 19672 33324 19700
rect 33318 19660 33324 19672
rect 33376 19660 33382 19712
rect 33502 19660 33508 19712
rect 33560 19700 33566 19712
rect 33689 19703 33747 19709
rect 33560 19672 33605 19700
rect 33560 19660 33566 19672
rect 33689 19669 33701 19703
rect 33735 19700 33747 19703
rect 33778 19700 33784 19712
rect 33735 19672 33784 19700
rect 33735 19669 33747 19672
rect 33689 19663 33747 19669
rect 33778 19660 33784 19672
rect 33836 19660 33842 19712
rect 34882 19660 34888 19712
rect 34940 19700 34946 19712
rect 37366 19700 37372 19712
rect 34940 19672 37372 19700
rect 34940 19660 34946 19672
rect 37366 19660 37372 19672
rect 37424 19660 37430 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 7098 19456 7104 19508
rect 7156 19496 7162 19508
rect 7745 19499 7803 19505
rect 7745 19496 7757 19499
rect 7156 19468 7757 19496
rect 7156 19456 7162 19468
rect 7745 19465 7757 19468
rect 7791 19465 7803 19499
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 7745 19459 7803 19465
rect 8864 19468 9413 19496
rect 8662 19428 8668 19440
rect 6380 19400 8668 19428
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 6380 19369 6408 19400
rect 8662 19388 8668 19400
rect 8720 19388 8726 19440
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 4672 19332 6377 19360
rect 4672 19320 4678 19332
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 6621 19363 6679 19369
rect 6621 19360 6633 19363
rect 6512 19332 6633 19360
rect 6512 19320 6518 19332
rect 6621 19329 6633 19332
rect 6667 19329 6679 19363
rect 6621 19323 6679 19329
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19360 8815 19363
rect 8864 19360 8892 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 9766 19496 9772 19508
rect 9727 19468 9772 19496
rect 9401 19459 9459 19465
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 10778 19496 10784 19508
rect 9916 19468 10784 19496
rect 9916 19456 9922 19468
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 10965 19499 11023 19505
rect 10965 19465 10977 19499
rect 11011 19496 11023 19499
rect 11011 19468 12756 19496
rect 11011 19465 11023 19468
rect 10965 19459 11023 19465
rect 8938 19388 8944 19440
rect 8996 19428 9002 19440
rect 12728 19437 12756 19468
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 13817 19499 13875 19505
rect 13817 19496 13829 19499
rect 13780 19468 13829 19496
rect 13780 19456 13786 19468
rect 13817 19465 13829 19468
rect 13863 19496 13875 19499
rect 14550 19496 14556 19508
rect 13863 19468 14556 19496
rect 13863 19465 13875 19468
rect 13817 19459 13875 19465
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14829 19499 14887 19505
rect 14829 19465 14841 19499
rect 14875 19496 14887 19499
rect 16758 19496 16764 19508
rect 14875 19468 16764 19496
rect 14875 19465 14887 19468
rect 14829 19459 14887 19465
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19496 16911 19499
rect 17034 19496 17040 19508
rect 16899 19468 17040 19496
rect 16899 19465 16911 19468
rect 16853 19459 16911 19465
rect 17034 19456 17040 19468
rect 17092 19496 17098 19508
rect 18322 19496 18328 19508
rect 17092 19468 18328 19496
rect 17092 19456 17098 19468
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 18509 19499 18567 19505
rect 18509 19465 18521 19499
rect 18555 19465 18567 19499
rect 18509 19459 18567 19465
rect 18877 19499 18935 19505
rect 18877 19465 18889 19499
rect 18923 19496 18935 19499
rect 20070 19496 20076 19508
rect 18923 19468 20076 19496
rect 18923 19465 18935 19468
rect 18877 19459 18935 19465
rect 12704 19431 12762 19437
rect 8996 19400 12572 19428
rect 8996 19388 9002 19400
rect 9030 19360 9036 19372
rect 8803 19332 8892 19360
rect 8956 19332 9036 19360
rect 8803 19329 8815 19332
rect 8757 19323 8815 19329
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 1854 19292 1860 19304
rect 1815 19264 1860 19292
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 2130 19292 2136 19304
rect 2091 19264 2136 19292
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 8956 19233 8984 19332
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19360 10839 19363
rect 11606 19360 11612 19372
rect 10827 19332 11612 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 10045 19295 10103 19301
rect 10045 19261 10057 19295
rect 10091 19292 10103 19295
rect 10318 19292 10324 19304
rect 10091 19264 10324 19292
rect 10091 19261 10103 19264
rect 10045 19255 10103 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12544 19292 12572 19400
rect 12704 19397 12716 19431
rect 12750 19397 12762 19431
rect 12704 19391 12762 19397
rect 15194 19388 15200 19440
rect 15252 19428 15258 19440
rect 15717 19431 15775 19437
rect 15717 19428 15729 19431
rect 15252 19400 15729 19428
rect 15252 19388 15258 19400
rect 15717 19397 15729 19400
rect 15763 19397 15775 19431
rect 15717 19391 15775 19397
rect 15933 19431 15991 19437
rect 15933 19397 15945 19431
rect 15979 19428 15991 19431
rect 16390 19428 16396 19440
rect 15979 19400 16396 19428
rect 15979 19397 15991 19400
rect 15933 19391 15991 19397
rect 16390 19388 16396 19400
rect 16448 19388 16454 19440
rect 18230 19428 18236 19440
rect 17052 19400 18236 19428
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14369 19363 14427 19369
rect 14369 19360 14381 19363
rect 14240 19332 14381 19360
rect 14240 19320 14246 19332
rect 14369 19329 14381 19332
rect 14415 19329 14427 19363
rect 14550 19360 14556 19372
rect 14511 19332 14556 19360
rect 14369 19323 14427 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 14826 19360 14832 19372
rect 14787 19332 14832 19360
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 15102 19360 15108 19372
rect 15063 19332 15108 19360
rect 15102 19320 15108 19332
rect 15160 19320 15166 19372
rect 17052 19369 17080 19400
rect 18230 19388 18236 19400
rect 18288 19388 18294 19440
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19329 17003 19363
rect 16945 19323 17003 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17218 19360 17224 19372
rect 17037 19323 17095 19329
rect 17144 19332 17224 19360
rect 12483 19264 12572 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 16669 19295 16727 19301
rect 16669 19292 16681 19295
rect 14700 19264 16681 19292
rect 14700 19252 14706 19264
rect 16669 19261 16681 19264
rect 16715 19261 16727 19295
rect 16960 19292 16988 19323
rect 17144 19292 17172 19332
rect 17218 19320 17224 19332
rect 17276 19360 17282 19372
rect 17865 19363 17923 19369
rect 17276 19332 17816 19360
rect 17276 19320 17282 19332
rect 16960 19264 17172 19292
rect 17788 19292 17816 19332
rect 17865 19329 17877 19363
rect 17911 19360 17923 19363
rect 18524 19360 18552 19459
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 25038 19496 25044 19508
rect 23492 19468 25044 19496
rect 19978 19437 19984 19440
rect 19972 19428 19984 19437
rect 19939 19400 19984 19428
rect 19972 19391 19984 19400
rect 19978 19388 19984 19391
rect 20036 19388 20042 19440
rect 22281 19431 22339 19437
rect 22281 19397 22293 19431
rect 22327 19428 22339 19431
rect 22462 19428 22468 19440
rect 22327 19400 22468 19428
rect 22327 19397 22339 19400
rect 22281 19391 22339 19397
rect 22462 19388 22468 19400
rect 22520 19428 22526 19440
rect 23014 19428 23020 19440
rect 22520 19400 23020 19428
rect 22520 19388 22526 19400
rect 23014 19388 23020 19400
rect 23072 19388 23078 19440
rect 17911 19332 18552 19360
rect 17911 19329 17923 19332
rect 17865 19323 17923 19329
rect 18966 19320 18972 19372
rect 19024 19360 19030 19372
rect 19024 19332 19069 19360
rect 19024 19320 19030 19332
rect 23382 19320 23388 19372
rect 23440 19360 23446 19372
rect 23492 19369 23520 19468
rect 25038 19456 25044 19468
rect 25096 19456 25102 19508
rect 26878 19456 26884 19508
rect 26936 19496 26942 19508
rect 26973 19499 27031 19505
rect 26973 19496 26985 19499
rect 26936 19468 26985 19496
rect 26936 19456 26942 19468
rect 26973 19465 26985 19468
rect 27019 19465 27031 19499
rect 27141 19499 27199 19505
rect 27141 19496 27153 19499
rect 26973 19459 27031 19465
rect 27080 19468 27153 19496
rect 26053 19431 26111 19437
rect 26053 19397 26065 19431
rect 26099 19428 26111 19431
rect 27080 19428 27108 19468
rect 27141 19465 27153 19468
rect 27187 19496 27199 19499
rect 27982 19496 27988 19508
rect 27187 19468 27988 19496
rect 27187 19465 27199 19468
rect 27141 19459 27199 19465
rect 27982 19456 27988 19468
rect 28040 19456 28046 19508
rect 28442 19456 28448 19508
rect 28500 19496 28506 19508
rect 28902 19496 28908 19508
rect 28500 19468 28908 19496
rect 28500 19456 28506 19468
rect 28902 19456 28908 19468
rect 28960 19456 28966 19508
rect 29638 19456 29644 19508
rect 29696 19496 29702 19508
rect 30374 19496 30380 19508
rect 29696 19468 30380 19496
rect 29696 19456 29702 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 31018 19456 31024 19508
rect 31076 19496 31082 19508
rect 32477 19499 32535 19505
rect 32477 19496 32489 19499
rect 31076 19468 32489 19496
rect 31076 19456 31082 19468
rect 32477 19465 32489 19468
rect 32523 19496 32535 19499
rect 33318 19496 33324 19508
rect 32523 19468 33324 19496
rect 32523 19465 32535 19468
rect 32477 19459 32535 19465
rect 33318 19456 33324 19468
rect 33376 19456 33382 19508
rect 33962 19456 33968 19508
rect 34020 19496 34026 19508
rect 34149 19499 34207 19505
rect 34149 19496 34161 19499
rect 34020 19468 34161 19496
rect 34020 19456 34026 19468
rect 34149 19465 34161 19468
rect 34195 19465 34207 19499
rect 36538 19496 36544 19508
rect 34149 19459 34207 19465
rect 34992 19468 36544 19496
rect 26099 19400 27108 19428
rect 27341 19431 27399 19437
rect 26099 19397 26111 19400
rect 26053 19391 26111 19397
rect 27341 19397 27353 19431
rect 27387 19397 27399 19431
rect 31573 19431 31631 19437
rect 27341 19391 27399 19397
rect 28966 19400 29500 19428
rect 23477 19363 23535 19369
rect 23477 19360 23489 19363
rect 23440 19332 23489 19360
rect 23440 19320 23446 19332
rect 23477 19329 23489 19332
rect 23523 19329 23535 19363
rect 23477 19323 23535 19329
rect 24854 19320 24860 19372
rect 24912 19320 24918 19372
rect 25406 19320 25412 19372
rect 25464 19360 25470 19372
rect 25961 19363 26019 19369
rect 25961 19360 25973 19363
rect 25464 19332 25973 19360
rect 25464 19320 25470 19332
rect 25961 19329 25973 19332
rect 26007 19329 26019 19363
rect 25961 19323 26019 19329
rect 26237 19363 26295 19369
rect 26237 19329 26249 19363
rect 26283 19329 26295 19363
rect 26237 19323 26295 19329
rect 18782 19292 18788 19304
rect 17788 19264 18788 19292
rect 16669 19255 16727 19261
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 19150 19292 19156 19304
rect 19111 19264 19156 19292
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19426 19252 19432 19304
rect 19484 19292 19490 19304
rect 19705 19295 19763 19301
rect 19705 19292 19717 19295
rect 19484 19264 19717 19292
rect 19484 19252 19490 19264
rect 19705 19261 19717 19264
rect 19751 19261 19763 19295
rect 19705 19255 19763 19261
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19292 22615 19295
rect 23014 19292 23020 19304
rect 22603 19264 23020 19292
rect 22603 19261 22615 19264
rect 22557 19255 22615 19261
rect 23014 19252 23020 19264
rect 23072 19252 23078 19304
rect 23750 19292 23756 19304
rect 23711 19264 23756 19292
rect 23750 19252 23756 19264
rect 23808 19252 23814 19304
rect 26050 19252 26056 19304
rect 26108 19292 26114 19304
rect 26252 19292 26280 19323
rect 26970 19320 26976 19372
rect 27028 19360 27034 19372
rect 27356 19360 27384 19391
rect 28258 19360 28264 19372
rect 27028 19332 27384 19360
rect 27448 19332 28264 19360
rect 27028 19320 27034 19332
rect 26108 19264 26280 19292
rect 26108 19252 26114 19264
rect 8941 19227 8999 19233
rect 8941 19193 8953 19227
rect 8987 19193 8999 19227
rect 8941 19187 8999 19193
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 11146 19224 11152 19236
rect 10284 19196 11152 19224
rect 10284 19184 10290 19196
rect 11146 19184 11152 19196
rect 11204 19224 11210 19236
rect 11701 19227 11759 19233
rect 11701 19224 11713 19227
rect 11204 19196 11713 19224
rect 11204 19184 11210 19196
rect 11701 19193 11713 19196
rect 11747 19193 11759 19227
rect 11701 19187 11759 19193
rect 13372 19196 15884 19224
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 11790 19156 11796 19168
rect 7892 19128 11796 19156
rect 7892 19116 7898 19128
rect 11790 19116 11796 19128
rect 11848 19156 11854 19168
rect 12802 19156 12808 19168
rect 11848 19128 12808 19156
rect 11848 19116 11854 19128
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 13372 19156 13400 19196
rect 15562 19156 15568 19168
rect 13136 19128 13400 19156
rect 15523 19128 15568 19156
rect 13136 19116 13142 19128
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 15746 19156 15752 19168
rect 15707 19128 15752 19156
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 15856 19156 15884 19196
rect 16022 19184 16028 19236
rect 16080 19224 16086 19236
rect 17221 19227 17279 19233
rect 17221 19224 17233 19227
rect 16080 19196 17233 19224
rect 16080 19184 16086 19196
rect 17221 19193 17233 19196
rect 17267 19193 17279 19227
rect 19242 19224 19248 19236
rect 17221 19187 17279 19193
rect 17328 19196 19248 19224
rect 17328 19156 17356 19196
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 24762 19184 24768 19236
rect 24820 19224 24826 19236
rect 25682 19224 25688 19236
rect 24820 19196 25688 19224
rect 24820 19184 24826 19196
rect 25682 19184 25688 19196
rect 25740 19184 25746 19236
rect 25866 19184 25872 19236
rect 25924 19224 25930 19236
rect 27448 19224 27476 19332
rect 28258 19320 28264 19332
rect 28316 19320 28322 19372
rect 28442 19360 28448 19372
rect 28403 19332 28448 19360
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28537 19363 28595 19369
rect 28537 19329 28549 19363
rect 28583 19360 28595 19363
rect 28966 19360 28994 19400
rect 28583 19332 28994 19360
rect 28583 19329 28595 19332
rect 28537 19323 28595 19329
rect 29178 19320 29184 19372
rect 29236 19360 29242 19372
rect 29472 19360 29500 19400
rect 31573 19397 31585 19431
rect 31619 19428 31631 19431
rect 32677 19431 32735 19437
rect 31619 19400 31754 19428
rect 31619 19397 31631 19400
rect 31573 19391 31631 19397
rect 29236 19332 29281 19360
rect 29380 19332 29500 19360
rect 29236 19320 29242 19332
rect 28074 19292 28080 19304
rect 28035 19264 28080 19292
rect 28074 19252 28080 19264
rect 28132 19252 28138 19304
rect 29086 19252 29092 19304
rect 29144 19292 29150 19304
rect 29380 19301 29408 19332
rect 29822 19320 29828 19372
rect 29880 19360 29886 19372
rect 30009 19363 30067 19369
rect 30009 19360 30021 19363
rect 29880 19332 30021 19360
rect 29880 19320 29886 19332
rect 30009 19329 30021 19332
rect 30055 19329 30067 19363
rect 30009 19323 30067 19329
rect 30098 19320 30104 19372
rect 30156 19360 30162 19372
rect 31297 19363 31355 19369
rect 31297 19360 31309 19363
rect 30156 19332 31309 19360
rect 30156 19320 30162 19332
rect 31297 19329 31309 19332
rect 31343 19329 31355 19363
rect 31726 19360 31754 19400
rect 32677 19397 32689 19431
rect 32723 19428 32735 19431
rect 32950 19428 32956 19440
rect 32723 19400 32956 19428
rect 32723 19397 32735 19400
rect 32677 19391 32735 19397
rect 32950 19388 32956 19400
rect 33008 19388 33014 19440
rect 34301 19431 34359 19437
rect 34301 19428 34313 19431
rect 33520 19400 34313 19428
rect 33134 19360 33140 19372
rect 31726 19332 33140 19360
rect 31297 19323 31355 19329
rect 33134 19320 33140 19332
rect 33192 19320 33198 19372
rect 33321 19363 33379 19369
rect 33321 19329 33333 19363
rect 33367 19360 33379 19363
rect 33410 19360 33416 19372
rect 33367 19332 33416 19360
rect 33367 19329 33379 19332
rect 33321 19323 33379 19329
rect 33410 19320 33416 19332
rect 33468 19320 33474 19372
rect 29273 19295 29331 19301
rect 29144 19264 29189 19292
rect 29144 19252 29150 19264
rect 29273 19261 29285 19295
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 29365 19295 29423 19301
rect 29365 19261 29377 19295
rect 29411 19292 29423 19295
rect 30285 19295 30343 19301
rect 30285 19292 30297 19295
rect 29411 19264 30297 19292
rect 29411 19261 29423 19264
rect 29365 19255 29423 19261
rect 30285 19261 30297 19264
rect 30331 19292 30343 19295
rect 30558 19292 30564 19304
rect 30331 19264 30564 19292
rect 30331 19261 30343 19264
rect 30285 19255 30343 19261
rect 25924 19196 26096 19224
rect 25924 19184 25930 19196
rect 18046 19156 18052 19168
rect 15856 19128 17356 19156
rect 18007 19128 18052 19156
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21085 19159 21143 19165
rect 21085 19156 21097 19159
rect 20956 19128 21097 19156
rect 20956 19116 20962 19128
rect 21085 19125 21097 19128
rect 21131 19156 21143 19159
rect 21726 19156 21732 19168
rect 21131 19128 21732 19156
rect 21131 19125 21143 19128
rect 21085 19119 21143 19125
rect 21726 19116 21732 19128
rect 21784 19116 21790 19168
rect 22002 19116 22008 19168
rect 22060 19156 22066 19168
rect 22554 19156 22560 19168
rect 22060 19128 22560 19156
rect 22060 19116 22066 19128
rect 22554 19116 22560 19128
rect 22612 19156 22618 19168
rect 23290 19156 23296 19168
rect 22612 19128 23296 19156
rect 22612 19116 22618 19128
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 25225 19159 25283 19165
rect 25225 19125 25237 19159
rect 25271 19156 25283 19159
rect 25406 19156 25412 19168
rect 25271 19128 25412 19156
rect 25271 19125 25283 19128
rect 25225 19119 25283 19125
rect 25406 19116 25412 19128
rect 25464 19116 25470 19168
rect 25958 19156 25964 19168
rect 25919 19128 25964 19156
rect 25958 19116 25964 19128
rect 26016 19116 26022 19168
rect 26068 19156 26096 19196
rect 26160 19196 27476 19224
rect 26160 19156 26188 19196
rect 28442 19184 28448 19236
rect 28500 19224 28506 19236
rect 29288 19224 29316 19255
rect 30558 19252 30564 19264
rect 30616 19292 30622 19304
rect 31478 19292 31484 19304
rect 30616 19264 31484 19292
rect 30616 19252 30622 19264
rect 31478 19252 31484 19264
rect 31536 19252 31542 19304
rect 31570 19252 31576 19304
rect 31628 19292 31634 19304
rect 31628 19264 31673 19292
rect 31628 19252 31634 19264
rect 32306 19252 32312 19304
rect 32364 19292 32370 19304
rect 33520 19301 33548 19400
rect 34301 19397 34313 19400
rect 34347 19428 34359 19431
rect 34514 19428 34520 19440
rect 34347 19397 34376 19428
rect 34475 19400 34520 19428
rect 34301 19391 34376 19397
rect 33505 19295 33563 19301
rect 33505 19292 33517 19295
rect 32364 19264 33517 19292
rect 32364 19252 32370 19264
rect 33505 19261 33517 19264
rect 33551 19261 33563 19295
rect 34348 19292 34376 19391
rect 34514 19388 34520 19400
rect 34572 19388 34578 19440
rect 34992 19369 35020 19468
rect 36538 19456 36544 19468
rect 36596 19456 36602 19508
rect 36722 19496 36728 19508
rect 36683 19468 36728 19496
rect 36722 19456 36728 19468
rect 36780 19496 36786 19508
rect 36780 19468 37320 19496
rect 36780 19456 36786 19468
rect 35894 19388 35900 19440
rect 35952 19388 35958 19440
rect 37292 19437 37320 19468
rect 37277 19431 37335 19437
rect 37277 19397 37289 19431
rect 37323 19397 37335 19431
rect 37277 19391 37335 19397
rect 37366 19388 37372 19440
rect 37424 19428 37430 19440
rect 37424 19400 37596 19428
rect 37424 19388 37430 19400
rect 34977 19363 35035 19369
rect 34977 19329 34989 19363
rect 35023 19329 35035 19363
rect 37458 19360 37464 19372
rect 34977 19323 35035 19329
rect 36464 19332 37228 19360
rect 37419 19332 37464 19360
rect 34514 19292 34520 19304
rect 34348 19264 34520 19292
rect 33505 19255 33563 19261
rect 34514 19252 34520 19264
rect 34572 19292 34578 19304
rect 34882 19292 34888 19304
rect 34572 19264 34888 19292
rect 34572 19252 34578 19264
rect 34882 19252 34888 19264
rect 34940 19252 34946 19304
rect 35253 19295 35311 19301
rect 35253 19261 35265 19295
rect 35299 19292 35311 19295
rect 35342 19292 35348 19304
rect 35299 19264 35348 19292
rect 35299 19261 35311 19264
rect 35253 19255 35311 19261
rect 35342 19252 35348 19264
rect 35400 19252 35406 19304
rect 35802 19252 35808 19304
rect 35860 19292 35866 19304
rect 36464 19292 36492 19332
rect 35860 19264 36492 19292
rect 37200 19292 37228 19332
rect 37458 19320 37464 19332
rect 37516 19320 37522 19372
rect 37568 19369 37596 19400
rect 37553 19363 37611 19369
rect 37553 19329 37565 19363
rect 37599 19329 37611 19363
rect 37553 19323 37611 19329
rect 37200 19264 37320 19292
rect 35860 19252 35866 19264
rect 28500 19196 29316 19224
rect 28500 19184 28506 19196
rect 30374 19184 30380 19236
rect 30432 19224 30438 19236
rect 37292 19233 37320 19264
rect 37277 19227 37335 19233
rect 30432 19196 35112 19224
rect 30432 19184 30438 19196
rect 26068 19128 26188 19156
rect 26510 19116 26516 19168
rect 26568 19156 26574 19168
rect 27157 19159 27215 19165
rect 27157 19156 27169 19159
rect 26568 19128 27169 19156
rect 26568 19116 26574 19128
rect 27157 19125 27169 19128
rect 27203 19125 27215 19159
rect 27157 19119 27215 19125
rect 29549 19159 29607 19165
rect 29549 19125 29561 19159
rect 29595 19156 29607 19159
rect 30190 19156 30196 19168
rect 29595 19128 30196 19156
rect 29595 19125 29607 19128
rect 29549 19119 29607 19125
rect 30190 19116 30196 19128
rect 30248 19116 30254 19168
rect 31389 19159 31447 19165
rect 31389 19125 31401 19159
rect 31435 19156 31447 19159
rect 32214 19156 32220 19168
rect 31435 19128 32220 19156
rect 31435 19125 31447 19128
rect 31389 19119 31447 19125
rect 32214 19116 32220 19128
rect 32272 19116 32278 19168
rect 32306 19116 32312 19168
rect 32364 19156 32370 19168
rect 32364 19128 32409 19156
rect 32364 19116 32370 19128
rect 32490 19116 32496 19168
rect 32548 19156 32554 19168
rect 33137 19159 33195 19165
rect 32548 19128 32593 19156
rect 32548 19116 32554 19128
rect 33137 19125 33149 19159
rect 33183 19156 33195 19159
rect 33226 19156 33232 19168
rect 33183 19128 33232 19156
rect 33183 19125 33195 19128
rect 33137 19119 33195 19125
rect 33226 19116 33232 19128
rect 33284 19116 33290 19168
rect 34333 19159 34391 19165
rect 34333 19125 34345 19159
rect 34379 19156 34391 19159
rect 34422 19156 34428 19168
rect 34379 19128 34428 19156
rect 34379 19125 34391 19128
rect 34333 19119 34391 19125
rect 34422 19116 34428 19128
rect 34480 19116 34486 19168
rect 35084 19156 35112 19196
rect 37277 19193 37289 19227
rect 37323 19193 37335 19227
rect 37277 19187 37335 19193
rect 35434 19156 35440 19168
rect 35084 19128 35440 19156
rect 35434 19116 35440 19128
rect 35492 19116 35498 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 1670 18952 1676 18964
rect 1627 18924 1676 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 1670 18912 1676 18924
rect 1728 18912 1734 18964
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 2133 18955 2191 18961
rect 2133 18952 2145 18955
rect 1912 18924 2145 18952
rect 1912 18912 1918 18924
rect 2133 18921 2145 18924
rect 2179 18921 2191 18955
rect 6454 18952 6460 18964
rect 6415 18924 6460 18952
rect 2133 18915 2191 18921
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18921 10563 18955
rect 10505 18915 10563 18921
rect 10689 18955 10747 18961
rect 10689 18921 10701 18955
rect 10735 18952 10747 18955
rect 14550 18952 14556 18964
rect 10735 18924 14556 18952
rect 10735 18921 10747 18924
rect 10689 18915 10747 18921
rect 10520 18884 10548 18915
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 15838 18912 15844 18964
rect 15896 18952 15902 18964
rect 16761 18955 16819 18961
rect 16761 18952 16773 18955
rect 15896 18924 16773 18952
rect 15896 18912 15902 18924
rect 10778 18884 10784 18896
rect 10520 18856 10784 18884
rect 10778 18844 10784 18856
rect 10836 18844 10842 18896
rect 13906 18884 13912 18896
rect 12406 18856 13912 18884
rect 9769 18819 9827 18825
rect 9769 18785 9781 18819
rect 9815 18816 9827 18819
rect 9858 18816 9864 18828
rect 9815 18788 9864 18816
rect 9815 18785 9827 18788
rect 9769 18779 9827 18785
rect 9858 18776 9864 18788
rect 9916 18776 9922 18828
rect 10318 18816 10324 18828
rect 10279 18788 10324 18816
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 11517 18819 11575 18825
rect 11517 18816 11529 18819
rect 10520 18788 11529 18816
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18748 2283 18751
rect 2314 18748 2320 18760
rect 2271 18720 2320 18748
rect 2271 18717 2283 18720
rect 2225 18711 2283 18717
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18748 6699 18751
rect 7466 18748 7472 18760
rect 6687 18720 7472 18748
rect 6687 18717 6699 18720
rect 6641 18711 6699 18717
rect 7466 18708 7472 18720
rect 7524 18708 7530 18760
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 9401 18751 9459 18757
rect 9401 18748 9413 18751
rect 8435 18720 9413 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 9401 18717 9413 18720
rect 9447 18717 9459 18751
rect 9582 18748 9588 18760
rect 9543 18720 9588 18748
rect 9401 18711 9459 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10520 18757 10548 18788
rect 11517 18785 11529 18788
rect 11563 18785 11575 18819
rect 11517 18779 11575 18785
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11940 18788 11989 18816
rect 11940 18776 11946 18788
rect 11977 18785 11989 18788
rect 12023 18816 12035 18819
rect 12406 18816 12434 18856
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 14921 18887 14979 18893
rect 14921 18853 14933 18887
rect 14967 18884 14979 18887
rect 15194 18884 15200 18896
rect 14967 18856 15200 18884
rect 14967 18853 14979 18856
rect 14921 18847 14979 18853
rect 15194 18844 15200 18856
rect 15252 18844 15258 18896
rect 16040 18825 16068 18924
rect 16761 18921 16773 18924
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 19429 18955 19487 18961
rect 19429 18921 19441 18955
rect 19475 18952 19487 18955
rect 20346 18952 20352 18964
rect 19475 18924 20352 18952
rect 19475 18921 19487 18924
rect 19429 18915 19487 18921
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 21821 18955 21879 18961
rect 21821 18952 21833 18955
rect 20456 18924 21833 18952
rect 17678 18844 17684 18896
rect 17736 18884 17742 18896
rect 18690 18884 18696 18896
rect 17736 18856 18696 18884
rect 17736 18844 17742 18856
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 18782 18844 18788 18896
rect 18840 18884 18846 18896
rect 20456 18884 20484 18924
rect 21821 18921 21833 18924
rect 21867 18921 21879 18955
rect 21821 18915 21879 18921
rect 22005 18955 22063 18961
rect 22005 18921 22017 18955
rect 22051 18921 22063 18955
rect 23658 18952 23664 18964
rect 22005 18915 22063 18921
rect 22756 18924 23664 18952
rect 18840 18856 20484 18884
rect 18840 18844 18846 18856
rect 21358 18844 21364 18896
rect 21416 18884 21422 18896
rect 22020 18884 22048 18915
rect 21416 18856 22048 18884
rect 21416 18844 21422 18856
rect 12023 18788 12434 18816
rect 16025 18819 16083 18825
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 16025 18785 16037 18819
rect 16071 18785 16083 18819
rect 16025 18779 16083 18785
rect 17218 18776 17224 18828
rect 17276 18816 17282 18828
rect 17494 18816 17500 18828
rect 17276 18788 17500 18816
rect 17276 18776 17282 18788
rect 17494 18776 17500 18788
rect 17552 18816 17558 18828
rect 17773 18819 17831 18825
rect 17773 18816 17785 18819
rect 17552 18788 17785 18816
rect 17552 18776 17558 18788
rect 17773 18785 17785 18788
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 17865 18819 17923 18825
rect 17865 18785 17877 18819
rect 17911 18816 17923 18819
rect 18230 18816 18236 18828
rect 17911 18788 18236 18816
rect 17911 18785 17923 18788
rect 17865 18779 17923 18785
rect 18230 18776 18236 18788
rect 18288 18816 18294 18828
rect 18506 18816 18512 18828
rect 18288 18788 18512 18816
rect 18288 18776 18294 18788
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 21542 18776 21548 18828
rect 21600 18816 21606 18828
rect 22756 18816 22784 18924
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 24210 18912 24216 18964
rect 24268 18952 24274 18964
rect 26234 18952 26240 18964
rect 24268 18924 26096 18952
rect 26195 18924 26240 18952
rect 24268 18912 24274 18924
rect 23382 18844 23388 18896
rect 23440 18844 23446 18896
rect 23569 18887 23627 18893
rect 23569 18853 23581 18887
rect 23615 18884 23627 18887
rect 25866 18884 25872 18896
rect 23615 18856 25872 18884
rect 23615 18853 23627 18856
rect 23569 18847 23627 18853
rect 25866 18844 25872 18856
rect 25924 18844 25930 18896
rect 26068 18884 26096 18924
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 27982 18952 27988 18964
rect 27943 18924 27988 18952
rect 27982 18912 27988 18924
rect 28040 18912 28046 18964
rect 28813 18955 28871 18961
rect 28813 18921 28825 18955
rect 28859 18921 28871 18955
rect 28813 18915 28871 18921
rect 28997 18955 29055 18961
rect 28997 18921 29009 18955
rect 29043 18952 29055 18955
rect 29270 18952 29276 18964
rect 29043 18924 29276 18952
rect 29043 18921 29055 18924
rect 28997 18915 29055 18921
rect 28534 18884 28540 18896
rect 26068 18856 28540 18884
rect 28534 18844 28540 18856
rect 28592 18844 28598 18896
rect 28828 18884 28856 18915
rect 29270 18912 29276 18924
rect 29328 18912 29334 18964
rect 30653 18955 30711 18961
rect 30208 18924 30420 18952
rect 30098 18884 30104 18896
rect 28828 18856 30104 18884
rect 30098 18844 30104 18856
rect 30156 18844 30162 18896
rect 23400 18816 23428 18844
rect 26326 18816 26332 18828
rect 21600 18788 22784 18816
rect 22848 18788 23428 18816
rect 25424 18788 25820 18816
rect 26287 18788 26332 18816
rect 21600 18776 21606 18788
rect 10505 18751 10563 18757
rect 10505 18748 10517 18751
rect 9732 18720 10517 18748
rect 9732 18708 9738 18720
rect 10505 18717 10517 18720
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 10686 18708 10692 18760
rect 10744 18748 10750 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 10744 18720 11345 18748
rect 10744 18708 10750 18720
rect 11333 18717 11345 18720
rect 11379 18748 11391 18751
rect 11790 18748 11796 18760
rect 11379 18720 11796 18748
rect 11379 18717 11391 18720
rect 11333 18711 11391 18717
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 12158 18748 12164 18760
rect 12119 18720 12164 18748
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 13078 18748 13084 18760
rect 12308 18720 12353 18748
rect 13039 18720 13084 18748
rect 12308 18708 12314 18720
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 13354 18748 13360 18760
rect 13315 18720 13360 18748
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15620 18720 15761 18748
rect 15620 18708 15626 18720
rect 15749 18717 15761 18720
rect 15795 18717 15807 18751
rect 15749 18711 15807 18717
rect 15856 18720 16712 18748
rect 10229 18683 10287 18689
rect 10229 18649 10241 18683
rect 10275 18680 10287 18683
rect 14737 18683 14795 18689
rect 10275 18652 10548 18680
rect 10275 18649 10287 18652
rect 10229 18643 10287 18649
rect 10520 18624 10548 18652
rect 14737 18649 14749 18683
rect 14783 18680 14795 18683
rect 15856 18680 15884 18720
rect 14783 18652 15884 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 16390 18640 16396 18692
rect 16448 18680 16454 18692
rect 16577 18683 16635 18689
rect 16577 18680 16589 18683
rect 16448 18652 16589 18680
rect 16448 18640 16454 18652
rect 16577 18649 16589 18652
rect 16623 18649 16635 18683
rect 16684 18680 16712 18720
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 17678 18748 17684 18760
rect 17092 18720 17684 18748
rect 17092 18708 17098 18720
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18748 18015 18751
rect 18598 18748 18604 18760
rect 18003 18720 18604 18748
rect 18003 18717 18015 18720
rect 17957 18711 18015 18717
rect 16793 18683 16851 18689
rect 16793 18680 16805 18683
rect 16684 18652 16805 18680
rect 16577 18643 16635 18649
rect 16793 18649 16805 18652
rect 16839 18680 16851 18683
rect 17310 18680 17316 18692
rect 16839 18652 17316 18680
rect 16839 18649 16851 18652
rect 16793 18643 16851 18649
rect 17310 18640 17316 18652
rect 17368 18640 17374 18692
rect 8205 18615 8263 18621
rect 8205 18581 8217 18615
rect 8251 18612 8263 18615
rect 8294 18612 8300 18624
rect 8251 18584 8300 18612
rect 8251 18581 8263 18584
rect 8205 18575 8263 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 10502 18572 10508 18624
rect 10560 18572 10566 18624
rect 10778 18572 10784 18624
rect 10836 18612 10842 18624
rect 11149 18615 11207 18621
rect 11149 18612 11161 18615
rect 10836 18584 11161 18612
rect 10836 18572 10842 18584
rect 11149 18581 11161 18584
rect 11195 18581 11207 18615
rect 11974 18612 11980 18624
rect 11935 18584 11980 18612
rect 11149 18575 11207 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12897 18615 12955 18621
rect 12897 18581 12909 18615
rect 12943 18612 12955 18615
rect 13170 18612 13176 18624
rect 12943 18584 13176 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 15378 18612 15384 18624
rect 13320 18584 13365 18612
rect 15339 18584 15384 18612
rect 13320 18572 13326 18584
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 15841 18615 15899 18621
rect 15841 18581 15853 18615
rect 15887 18612 15899 18615
rect 16482 18612 16488 18624
rect 15887 18584 16488 18612
rect 15887 18581 15899 18584
rect 15841 18575 15899 18581
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 16942 18572 16948 18624
rect 17000 18612 17006 18624
rect 17972 18612 18000 18711
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18748 19579 18751
rect 20806 18748 20812 18760
rect 19567 18720 20812 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 21361 18751 21419 18757
rect 21361 18717 21373 18751
rect 21407 18748 21419 18751
rect 22094 18748 22100 18760
rect 21407 18720 22100 18748
rect 21407 18717 21419 18720
rect 21361 18711 21419 18717
rect 22094 18708 22100 18720
rect 22152 18748 22158 18760
rect 22848 18748 22876 18788
rect 25424 18760 25452 18788
rect 22152 18720 22876 18748
rect 22152 18708 22158 18720
rect 22922 18708 22928 18760
rect 22980 18748 22986 18760
rect 22980 18720 23025 18748
rect 22980 18708 22986 18720
rect 23290 18708 23296 18760
rect 23348 18748 23354 18760
rect 23385 18751 23443 18757
rect 23385 18748 23397 18751
rect 23348 18720 23397 18748
rect 23348 18708 23354 18720
rect 23385 18717 23397 18720
rect 23431 18717 23443 18751
rect 25406 18748 25412 18760
rect 25367 18720 25412 18748
rect 23385 18711 23443 18717
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 25685 18751 25743 18757
rect 25685 18717 25697 18751
rect 25731 18717 25743 18751
rect 25792 18748 25820 18788
rect 26326 18776 26332 18788
rect 26384 18776 26390 18828
rect 27341 18819 27399 18825
rect 27341 18785 27353 18819
rect 27387 18816 27399 18819
rect 30208 18816 30236 18924
rect 30282 18844 30288 18896
rect 30340 18844 30346 18896
rect 27387 18788 30236 18816
rect 27387 18785 27399 18788
rect 27341 18779 27399 18785
rect 26421 18751 26479 18757
rect 26421 18748 26433 18751
rect 25792 18720 26433 18748
rect 25685 18711 25743 18717
rect 26421 18717 26433 18720
rect 26467 18717 26479 18751
rect 26421 18711 26479 18717
rect 18046 18640 18052 18692
rect 18104 18680 18110 18692
rect 21094 18683 21152 18689
rect 21094 18680 21106 18683
rect 18104 18652 21106 18680
rect 18104 18640 18110 18652
rect 21094 18649 21106 18652
rect 21140 18649 21152 18683
rect 21094 18643 21152 18649
rect 21726 18640 21732 18692
rect 21784 18680 21790 18692
rect 21973 18683 22031 18689
rect 21973 18680 21985 18683
rect 21784 18652 21985 18680
rect 21784 18640 21790 18652
rect 21973 18649 21985 18652
rect 22019 18649 22031 18683
rect 21973 18643 22031 18649
rect 22189 18683 22247 18689
rect 22189 18649 22201 18683
rect 22235 18649 22247 18683
rect 22940 18680 22968 18708
rect 24489 18683 24547 18689
rect 24489 18680 24501 18683
rect 22940 18652 24501 18680
rect 22189 18643 22247 18649
rect 24489 18649 24501 18652
rect 24535 18649 24547 18683
rect 25700 18680 25728 18711
rect 26878 18708 26884 18760
rect 26936 18748 26942 18760
rect 27433 18751 27491 18757
rect 26936 18720 27384 18748
rect 26936 18708 26942 18720
rect 26050 18680 26056 18692
rect 25700 18652 26056 18680
rect 24489 18643 24547 18649
rect 17000 18584 18000 18612
rect 18141 18615 18199 18621
rect 17000 18572 17006 18584
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18506 18612 18512 18624
rect 18187 18584 18512 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 19150 18572 19156 18624
rect 19208 18612 19214 18624
rect 19981 18615 20039 18621
rect 19981 18612 19993 18615
rect 19208 18584 19993 18612
rect 19208 18572 19214 18584
rect 19981 18581 19993 18584
rect 20027 18612 20039 18615
rect 22204 18612 22232 18643
rect 26050 18640 26056 18652
rect 26108 18640 26114 18692
rect 26142 18640 26148 18692
rect 26200 18680 26206 18692
rect 26970 18680 26976 18692
rect 26200 18652 26245 18680
rect 26528 18652 26976 18680
rect 26200 18640 26206 18652
rect 22738 18612 22744 18624
rect 20027 18584 22232 18612
rect 22699 18584 22744 18612
rect 20027 18581 20039 18584
rect 19981 18575 20039 18581
rect 22738 18572 22744 18584
rect 22796 18572 22802 18624
rect 24578 18612 24584 18624
rect 24539 18584 24584 18612
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 25222 18612 25228 18624
rect 25183 18584 25228 18612
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 25593 18615 25651 18621
rect 25593 18581 25605 18615
rect 25639 18612 25651 18615
rect 26528 18612 26556 18652
rect 26970 18640 26976 18652
rect 27028 18640 27034 18692
rect 27356 18680 27384 18720
rect 27433 18717 27445 18751
rect 27479 18748 27491 18751
rect 29086 18748 29092 18760
rect 27479 18720 29092 18748
rect 27479 18717 27491 18720
rect 27433 18711 27491 18717
rect 29086 18708 29092 18720
rect 29144 18748 29150 18760
rect 29144 18720 29960 18748
rect 29144 18708 29150 18720
rect 28077 18683 28135 18689
rect 27356 18652 28028 18680
rect 25639 18584 26556 18612
rect 26605 18615 26663 18621
rect 25639 18581 25651 18584
rect 25593 18575 25651 18581
rect 26605 18581 26617 18615
rect 26651 18612 26663 18615
rect 27614 18612 27620 18624
rect 26651 18584 27620 18612
rect 26651 18581 26663 18584
rect 26605 18575 26663 18581
rect 27614 18572 27620 18584
rect 27672 18572 27678 18624
rect 28000 18612 28028 18652
rect 28077 18649 28089 18683
rect 28123 18680 28135 18683
rect 28258 18680 28264 18692
rect 28123 18652 28264 18680
rect 28123 18649 28135 18652
rect 28077 18643 28135 18649
rect 28258 18640 28264 18652
rect 28316 18640 28322 18692
rect 28629 18683 28687 18689
rect 28629 18649 28641 18683
rect 28675 18649 28687 18683
rect 28629 18643 28687 18649
rect 28845 18683 28903 18689
rect 28845 18649 28857 18683
rect 28891 18680 28903 18683
rect 29546 18680 29552 18692
rect 28891 18652 29552 18680
rect 28891 18649 28903 18652
rect 28845 18643 28903 18649
rect 28644 18612 28672 18643
rect 29546 18640 29552 18652
rect 29604 18640 29610 18692
rect 29932 18680 29960 18720
rect 30006 18708 30012 18760
rect 30064 18748 30070 18760
rect 30190 18748 30196 18760
rect 30064 18720 30109 18748
rect 30151 18720 30196 18748
rect 30064 18708 30070 18720
rect 30190 18708 30196 18720
rect 30248 18708 30254 18760
rect 30300 18757 30328 18844
rect 30392 18757 30420 18924
rect 30653 18921 30665 18955
rect 30699 18952 30711 18955
rect 30742 18952 30748 18964
rect 30699 18924 30748 18952
rect 30699 18921 30711 18924
rect 30653 18915 30711 18921
rect 30742 18912 30748 18924
rect 30800 18912 30806 18964
rect 30834 18912 30840 18964
rect 30892 18952 30898 18964
rect 31297 18955 31355 18961
rect 31297 18952 31309 18955
rect 30892 18924 31309 18952
rect 30892 18912 30898 18924
rect 31297 18921 31309 18924
rect 31343 18921 31355 18955
rect 31297 18915 31355 18921
rect 31386 18912 31392 18964
rect 31444 18952 31450 18964
rect 31570 18952 31576 18964
rect 31444 18924 31576 18952
rect 31444 18912 31450 18924
rect 31570 18912 31576 18924
rect 31628 18952 31634 18964
rect 34330 18952 34336 18964
rect 31628 18924 34336 18952
rect 31628 18912 31634 18924
rect 34330 18912 34336 18924
rect 34388 18912 34394 18964
rect 34885 18955 34943 18961
rect 34885 18921 34897 18955
rect 34931 18952 34943 18955
rect 35621 18955 35679 18961
rect 34931 18924 35572 18952
rect 34931 18921 34943 18924
rect 34885 18915 34943 18921
rect 30285 18751 30343 18757
rect 30285 18717 30297 18751
rect 30331 18717 30343 18751
rect 30285 18711 30343 18717
rect 30377 18751 30435 18757
rect 30377 18717 30389 18751
rect 30423 18717 30435 18751
rect 30377 18711 30435 18717
rect 30852 18680 30880 18912
rect 35544 18896 35572 18924
rect 35621 18921 35633 18955
rect 35667 18952 35679 18955
rect 35894 18952 35900 18964
rect 35667 18924 35900 18952
rect 35667 18921 35679 18924
rect 35621 18915 35679 18921
rect 35894 18912 35900 18924
rect 35952 18912 35958 18964
rect 31202 18844 31208 18896
rect 31260 18884 31266 18896
rect 31260 18856 34836 18884
rect 31260 18844 31266 18856
rect 34808 18816 34836 18856
rect 35526 18844 35532 18896
rect 35584 18844 35590 18896
rect 36538 18844 36544 18896
rect 36596 18844 36602 18896
rect 35894 18816 35900 18828
rect 34808 18788 35900 18816
rect 35894 18776 35900 18788
rect 35952 18776 35958 18828
rect 36556 18816 36584 18844
rect 37921 18819 37979 18825
rect 37921 18816 37933 18819
rect 36556 18788 37933 18816
rect 37921 18785 37933 18788
rect 37967 18785 37979 18819
rect 37921 18779 37979 18785
rect 31110 18708 31116 18760
rect 31168 18748 31174 18760
rect 31168 18720 31524 18748
rect 31168 18708 31174 18720
rect 29932 18652 30880 18680
rect 31018 18640 31024 18692
rect 31076 18680 31082 18692
rect 31496 18689 31524 18720
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32309 18751 32367 18757
rect 32309 18748 32321 18751
rect 32272 18720 32321 18748
rect 32272 18708 32278 18720
rect 32309 18717 32321 18720
rect 32355 18717 32367 18751
rect 32309 18711 32367 18717
rect 32585 18751 32643 18757
rect 32585 18717 32597 18751
rect 32631 18748 32643 18751
rect 33042 18748 33048 18760
rect 32631 18720 33048 18748
rect 32631 18717 32643 18720
rect 32585 18711 32643 18717
rect 31265 18683 31323 18689
rect 31265 18680 31277 18683
rect 31076 18652 31277 18680
rect 31076 18640 31082 18652
rect 31265 18649 31277 18652
rect 31311 18649 31323 18683
rect 31265 18643 31323 18649
rect 31481 18683 31539 18689
rect 31481 18649 31493 18683
rect 31527 18649 31539 18683
rect 32324 18680 32352 18711
rect 33042 18708 33048 18720
rect 33100 18748 33106 18760
rect 33505 18751 33563 18757
rect 33505 18748 33517 18751
rect 33100 18720 33517 18748
rect 33100 18708 33106 18720
rect 33505 18717 33517 18720
rect 33551 18748 33563 18751
rect 34149 18751 34207 18757
rect 33551 18720 34008 18748
rect 33551 18717 33563 18720
rect 33505 18711 33563 18717
rect 32490 18680 32496 18692
rect 32324 18652 32496 18680
rect 31481 18643 31539 18649
rect 32490 18640 32496 18652
rect 32548 18680 32554 18692
rect 33226 18680 33232 18692
rect 32548 18652 33232 18680
rect 32548 18640 32554 18652
rect 33226 18640 33232 18652
rect 33284 18640 33290 18692
rect 33318 18640 33324 18692
rect 33376 18680 33382 18692
rect 33413 18683 33471 18689
rect 33413 18680 33425 18683
rect 33376 18652 33425 18680
rect 33376 18640 33382 18652
rect 33413 18649 33425 18652
rect 33459 18649 33471 18683
rect 33413 18643 33471 18649
rect 28000 18584 28672 18612
rect 28994 18572 29000 18624
rect 29052 18612 29058 18624
rect 30006 18612 30012 18624
rect 29052 18584 30012 18612
rect 29052 18572 29058 18584
rect 30006 18572 30012 18584
rect 30064 18572 30070 18624
rect 31110 18612 31116 18624
rect 31071 18584 31116 18612
rect 31110 18572 31116 18584
rect 31168 18572 31174 18624
rect 32398 18612 32404 18624
rect 32359 18584 32404 18612
rect 32398 18572 32404 18584
rect 32456 18572 32462 18624
rect 32769 18615 32827 18621
rect 32769 18581 32781 18615
rect 32815 18612 32827 18615
rect 33134 18612 33140 18624
rect 32815 18584 33140 18612
rect 32815 18581 32827 18584
rect 32769 18575 32827 18581
rect 33134 18572 33140 18584
rect 33192 18572 33198 18624
rect 33505 18615 33563 18621
rect 33505 18581 33517 18615
rect 33551 18612 33563 18615
rect 33686 18612 33692 18624
rect 33551 18584 33692 18612
rect 33551 18581 33563 18584
rect 33505 18575 33563 18581
rect 33686 18572 33692 18584
rect 33744 18572 33750 18624
rect 33980 18621 34008 18720
rect 34149 18717 34161 18751
rect 34195 18748 34207 18751
rect 34790 18748 34796 18760
rect 34195 18720 34796 18748
rect 34195 18717 34207 18720
rect 34149 18711 34207 18717
rect 34790 18708 34796 18720
rect 34848 18708 34854 18760
rect 35529 18751 35587 18757
rect 35529 18717 35541 18751
rect 35575 18748 35587 18751
rect 35618 18748 35624 18760
rect 35575 18720 35624 18748
rect 35575 18717 35587 18720
rect 35529 18711 35587 18717
rect 35618 18708 35624 18720
rect 35676 18748 35682 18760
rect 35986 18748 35992 18760
rect 35676 18720 35992 18748
rect 35676 18708 35682 18720
rect 35986 18708 35992 18720
rect 36044 18708 36050 18760
rect 34422 18640 34428 18692
rect 34480 18680 34486 18692
rect 34701 18683 34759 18689
rect 34701 18680 34713 18683
rect 34480 18652 34713 18680
rect 34480 18640 34486 18652
rect 34701 18649 34713 18652
rect 34747 18649 34759 18683
rect 34808 18680 34836 18708
rect 34808 18652 36216 18680
rect 34701 18643 34759 18649
rect 33965 18615 34023 18621
rect 33965 18581 33977 18615
rect 34011 18581 34023 18615
rect 34716 18612 34744 18643
rect 34790 18612 34796 18624
rect 34716 18584 34796 18612
rect 33965 18575 34023 18581
rect 34790 18572 34796 18584
rect 34848 18572 34854 18624
rect 34882 18572 34888 18624
rect 34940 18621 34946 18624
rect 34940 18615 34959 18621
rect 34947 18581 34959 18615
rect 34940 18575 34959 18581
rect 35069 18615 35127 18621
rect 35069 18581 35081 18615
rect 35115 18612 35127 18615
rect 35434 18612 35440 18624
rect 35115 18584 35440 18612
rect 35115 18581 35127 18584
rect 35069 18575 35127 18581
rect 34940 18572 34946 18575
rect 35434 18572 35440 18584
rect 35492 18572 35498 18624
rect 36188 18621 36216 18652
rect 36354 18640 36360 18692
rect 36412 18680 36418 18692
rect 37642 18680 37648 18692
rect 36412 18652 36478 18680
rect 37603 18652 37648 18680
rect 36412 18640 36418 18652
rect 37642 18640 37648 18652
rect 37700 18640 37706 18692
rect 36173 18615 36231 18621
rect 36173 18581 36185 18615
rect 36219 18581 36231 18615
rect 36173 18575 36231 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 10321 18411 10379 18417
rect 10321 18408 10333 18411
rect 9640 18380 10333 18408
rect 9640 18368 9646 18380
rect 10321 18377 10333 18380
rect 10367 18377 10379 18411
rect 10778 18408 10784 18420
rect 10739 18380 10784 18408
rect 10321 18371 10379 18377
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 11606 18368 11612 18420
rect 11664 18408 11670 18420
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 11664 18380 12909 18408
rect 11664 18368 11670 18380
rect 12897 18377 12909 18380
rect 12943 18377 12955 18411
rect 12897 18371 12955 18377
rect 16853 18411 16911 18417
rect 16853 18377 16865 18411
rect 16899 18408 16911 18411
rect 16942 18408 16948 18420
rect 16899 18380 16948 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 19981 18411 20039 18417
rect 19981 18377 19993 18411
rect 20027 18408 20039 18411
rect 20070 18408 20076 18420
rect 20027 18380 20076 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 21177 18411 21235 18417
rect 21177 18377 21189 18411
rect 21223 18408 21235 18411
rect 21542 18408 21548 18420
rect 21223 18380 21548 18408
rect 21223 18377 21235 18380
rect 21177 18371 21235 18377
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 24946 18408 24952 18420
rect 24907 18380 24952 18408
rect 24946 18368 24952 18380
rect 25004 18368 25010 18420
rect 25958 18417 25964 18420
rect 25945 18411 25964 18417
rect 25945 18377 25957 18411
rect 25945 18371 25964 18377
rect 25958 18368 25964 18371
rect 26016 18368 26022 18420
rect 26418 18408 26424 18420
rect 26068 18380 26424 18408
rect 8662 18340 8668 18352
rect 8036 18312 8668 18340
rect 8036 18281 8064 18312
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 10873 18343 10931 18349
rect 10873 18309 10885 18343
rect 10919 18340 10931 18343
rect 13262 18340 13268 18352
rect 10919 18312 13268 18340
rect 10919 18309 10931 18312
rect 10873 18303 10931 18309
rect 13262 18300 13268 18312
rect 13320 18340 13326 18352
rect 13446 18340 13452 18352
rect 13320 18312 13452 18340
rect 13320 18300 13326 18312
rect 13446 18300 13452 18312
rect 13504 18340 13510 18352
rect 13504 18312 14044 18340
rect 13504 18300 13510 18312
rect 8294 18281 8300 18284
rect 8021 18275 8079 18281
rect 8021 18241 8033 18275
rect 8067 18241 8079 18275
rect 8288 18272 8300 18281
rect 8255 18244 8300 18272
rect 8021 18235 8079 18241
rect 8288 18235 8300 18244
rect 8294 18232 8300 18235
rect 8352 18232 8358 18284
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 11606 18272 11612 18284
rect 10643 18244 11612 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 11606 18232 11612 18244
rect 11664 18272 11670 18284
rect 11885 18275 11943 18281
rect 11885 18272 11897 18275
rect 11664 18244 11897 18272
rect 11664 18232 11670 18244
rect 11885 18241 11897 18244
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 13814 18272 13820 18284
rect 13127 18244 13820 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 14016 18281 14044 18312
rect 19334 18300 19340 18352
rect 19392 18340 19398 18352
rect 21358 18340 21364 18352
rect 19392 18312 20208 18340
rect 19392 18300 19398 18312
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 15013 18275 15071 18281
rect 15013 18272 15025 18275
rect 14047 18244 15025 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 15013 18241 15025 18244
rect 15059 18272 15071 18275
rect 15746 18272 15752 18284
rect 15059 18244 15752 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 19242 18272 19248 18284
rect 19300 18281 19306 18284
rect 19212 18244 19248 18272
rect 19242 18232 19248 18244
rect 19300 18235 19312 18281
rect 19300 18232 19306 18235
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 20180 18281 20208 18312
rect 20364 18312 21364 18340
rect 20364 18284 20392 18312
rect 21358 18300 21364 18312
rect 21416 18300 21422 18352
rect 22094 18340 22100 18352
rect 21836 18312 22100 18340
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19484 18244 19533 18272
rect 19484 18232 19490 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 20165 18275 20223 18281
rect 20165 18241 20177 18275
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20346 18232 20352 18284
rect 20404 18272 20410 18284
rect 21836 18281 21864 18312
rect 22094 18300 22100 18312
rect 22152 18300 22158 18352
rect 22554 18300 22560 18352
rect 22612 18300 22618 18352
rect 23842 18340 23848 18352
rect 23400 18312 23848 18340
rect 21269 18275 21327 18281
rect 20404 18244 20497 18272
rect 20404 18232 20410 18244
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 21821 18275 21879 18281
rect 21821 18241 21833 18275
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 10502 18204 10508 18216
rect 9416 18176 10508 18204
rect 9416 18145 9444 18176
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 9401 18139 9459 18145
rect 9401 18105 9413 18139
rect 9447 18105 9459 18139
rect 10980 18136 11008 18167
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11296 18176 11713 18204
rect 11296 18164 11302 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 11790 18164 11796 18216
rect 11848 18204 11854 18216
rect 11977 18207 12035 18213
rect 11848 18176 11893 18204
rect 11848 18164 11854 18176
rect 11977 18173 11989 18207
rect 12023 18204 12035 18207
rect 12250 18204 12256 18216
rect 12023 18176 12256 18204
rect 12023 18173 12035 18176
rect 11977 18167 12035 18173
rect 12250 18164 12256 18176
rect 12308 18204 12314 18216
rect 13262 18204 13268 18216
rect 12308 18176 12434 18204
rect 13223 18176 13268 18204
rect 12308 18164 12314 18176
rect 12158 18136 12164 18148
rect 10980 18108 12164 18136
rect 9401 18099 9459 18105
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 11480 18040 11529 18068
rect 11480 18028 11486 18040
rect 11517 18037 11529 18040
rect 11563 18037 11575 18071
rect 12406 18068 12434 18176
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 13964 18176 14749 18204
rect 13964 18164 13970 18176
rect 14737 18173 14749 18176
rect 14783 18204 14795 18207
rect 14918 18204 14924 18216
rect 14783 18176 14924 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 17034 18204 17040 18216
rect 16632 18176 17040 18204
rect 16632 18164 16638 18176
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 12802 18096 12808 18148
rect 12860 18136 12866 18148
rect 14185 18139 14243 18145
rect 14185 18136 14197 18139
rect 12860 18108 14197 18136
rect 12860 18096 12866 18108
rect 14185 18105 14197 18108
rect 14231 18136 14243 18139
rect 17218 18136 17224 18148
rect 14231 18108 16896 18136
rect 17179 18108 17224 18136
rect 14231 18105 14243 18108
rect 14185 18099 14243 18105
rect 16868 18080 16896 18108
rect 17218 18096 17224 18108
rect 17276 18096 17282 18148
rect 16574 18068 16580 18080
rect 12406 18040 16580 18068
rect 11517 18031 11575 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 16669 18071 16727 18077
rect 16669 18037 16681 18071
rect 16715 18068 16727 18071
rect 16758 18068 16764 18080
rect 16715 18040 16764 18068
rect 16715 18037 16727 18040
rect 16669 18031 16727 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 16850 18028 16856 18080
rect 16908 18068 16914 18080
rect 18141 18071 18199 18077
rect 16908 18040 16953 18068
rect 16908 18028 16914 18040
rect 18141 18037 18153 18071
rect 18187 18068 18199 18071
rect 18230 18068 18236 18080
rect 18187 18040 18236 18068
rect 18187 18037 18199 18040
rect 18141 18031 18199 18037
rect 18230 18028 18236 18040
rect 18288 18068 18294 18080
rect 20346 18068 20352 18080
rect 18288 18040 20352 18068
rect 18288 18028 18294 18040
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 21284 18068 21312 18235
rect 22097 18207 22155 18213
rect 22097 18173 22109 18207
rect 22143 18204 22155 18207
rect 23400 18204 23428 18312
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 24578 18340 24584 18352
rect 24320 18312 24584 18340
rect 24210 18272 24216 18284
rect 22143 18176 23428 18204
rect 23492 18244 24216 18272
rect 22143 18173 22155 18176
rect 22097 18167 22155 18173
rect 23492 18068 23520 18244
rect 24210 18232 24216 18244
rect 24268 18232 24274 18284
rect 24320 18281 24348 18312
rect 24578 18300 24584 18312
rect 24636 18340 24642 18352
rect 26068 18340 26096 18380
rect 26418 18368 26424 18380
rect 26476 18368 26482 18420
rect 27062 18368 27068 18420
rect 27120 18408 27126 18420
rect 29089 18411 29147 18417
rect 29089 18408 29101 18411
rect 27120 18380 29101 18408
rect 27120 18368 27126 18380
rect 29089 18377 29101 18380
rect 29135 18408 29147 18411
rect 31018 18408 31024 18420
rect 29135 18380 31024 18408
rect 29135 18377 29147 18380
rect 29089 18371 29147 18377
rect 31018 18368 31024 18380
rect 31076 18368 31082 18420
rect 31481 18411 31539 18417
rect 31481 18377 31493 18411
rect 31527 18408 31539 18411
rect 31662 18408 31668 18420
rect 31527 18380 31668 18408
rect 31527 18377 31539 18380
rect 31481 18371 31539 18377
rect 31662 18368 31668 18380
rect 31720 18368 31726 18420
rect 32950 18368 32956 18420
rect 33008 18408 33014 18420
rect 33045 18411 33103 18417
rect 33045 18408 33057 18411
rect 33008 18380 33057 18408
rect 33008 18368 33014 18380
rect 33045 18377 33057 18380
rect 33091 18377 33103 18411
rect 33045 18371 33103 18377
rect 33229 18411 33287 18417
rect 33229 18377 33241 18411
rect 33275 18408 33287 18411
rect 33502 18408 33508 18420
rect 33275 18380 33508 18408
rect 33275 18377 33287 18380
rect 33229 18371 33287 18377
rect 33502 18368 33508 18380
rect 33560 18368 33566 18420
rect 34790 18368 34796 18420
rect 34848 18408 34854 18420
rect 36722 18408 36728 18420
rect 34848 18380 36728 18408
rect 34848 18368 34854 18380
rect 36722 18368 36728 18380
rect 36780 18368 36786 18420
rect 37461 18411 37519 18417
rect 37461 18377 37473 18411
rect 37507 18408 37519 18411
rect 37642 18408 37648 18420
rect 37507 18380 37648 18408
rect 37507 18377 37519 18380
rect 37461 18371 37519 18377
rect 37642 18368 37648 18380
rect 37700 18368 37706 18420
rect 24636 18312 26096 18340
rect 24636 18300 24642 18312
rect 26142 18300 26148 18352
rect 26200 18340 26206 18352
rect 26878 18340 26884 18352
rect 26200 18312 26884 18340
rect 26200 18300 26206 18312
rect 26878 18300 26884 18312
rect 26936 18300 26942 18352
rect 26973 18343 27031 18349
rect 26973 18309 26985 18343
rect 27019 18309 27031 18343
rect 30650 18340 30656 18352
rect 26973 18303 27031 18309
rect 30116 18312 30656 18340
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 25133 18275 25191 18281
rect 25133 18241 25145 18275
rect 25179 18241 25191 18275
rect 25133 18235 25191 18241
rect 25317 18275 25375 18281
rect 25317 18241 25329 18275
rect 25363 18272 25375 18275
rect 26988 18272 27016 18303
rect 27246 18272 27252 18284
rect 25363 18244 27016 18272
rect 27207 18244 27252 18272
rect 25363 18241 25375 18244
rect 25317 18235 25375 18241
rect 25148 18204 25176 18235
rect 27246 18232 27252 18244
rect 27304 18232 27310 18284
rect 28258 18272 28264 18284
rect 28219 18244 28264 18272
rect 28258 18232 28264 18244
rect 28316 18272 28322 18284
rect 28997 18275 29055 18281
rect 28997 18272 29009 18275
rect 28316 18244 29009 18272
rect 28316 18232 28322 18244
rect 28997 18241 29009 18244
rect 29043 18272 29055 18275
rect 29825 18275 29883 18281
rect 29825 18272 29837 18275
rect 29043 18244 29837 18272
rect 29043 18241 29055 18244
rect 28997 18235 29055 18241
rect 29825 18241 29837 18244
rect 29871 18241 29883 18275
rect 29825 18235 29883 18241
rect 30116 18216 30144 18312
rect 30650 18300 30656 18312
rect 30708 18340 30714 18352
rect 31113 18343 31171 18349
rect 31113 18340 31125 18343
rect 30708 18312 31125 18340
rect 30708 18300 30714 18312
rect 31113 18309 31125 18312
rect 31159 18309 31171 18343
rect 31113 18303 31171 18309
rect 31329 18343 31387 18349
rect 31329 18309 31341 18343
rect 31375 18340 31387 18343
rect 31375 18312 31524 18340
rect 31375 18309 31387 18312
rect 31329 18303 31387 18309
rect 31496 18284 31524 18312
rect 35894 18300 35900 18352
rect 35952 18340 35958 18352
rect 35952 18312 37964 18340
rect 35952 18300 35958 18312
rect 31478 18232 31484 18284
rect 31536 18232 31542 18284
rect 32858 18272 32864 18284
rect 32819 18244 32864 18272
rect 32858 18232 32864 18244
rect 32916 18232 32922 18284
rect 32953 18275 33011 18281
rect 32953 18241 32965 18275
rect 32999 18272 33011 18275
rect 33042 18272 33048 18284
rect 32999 18244 33048 18272
rect 32999 18241 33011 18244
rect 32953 18235 33011 18241
rect 33042 18232 33048 18244
rect 33100 18232 33106 18284
rect 36078 18272 36084 18284
rect 35650 18244 36084 18272
rect 36078 18232 36084 18244
rect 36136 18232 36142 18284
rect 36170 18232 36176 18284
rect 36228 18272 36234 18284
rect 37936 18281 37964 18312
rect 36449 18275 36507 18281
rect 36449 18272 36461 18275
rect 36228 18244 36461 18272
rect 36228 18232 36234 18244
rect 36449 18241 36461 18244
rect 36495 18241 36507 18275
rect 36449 18235 36507 18241
rect 37277 18275 37335 18281
rect 37277 18241 37289 18275
rect 37323 18241 37335 18275
rect 37277 18235 37335 18241
rect 37921 18275 37979 18281
rect 37921 18241 37933 18275
rect 37967 18241 37979 18275
rect 37921 18235 37979 18241
rect 26326 18204 26332 18216
rect 25148 18176 26332 18204
rect 26326 18164 26332 18176
rect 26384 18164 26390 18216
rect 26973 18207 27031 18213
rect 26973 18173 26985 18207
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 23569 18139 23627 18145
rect 23569 18105 23581 18139
rect 23615 18136 23627 18139
rect 25130 18136 25136 18148
rect 23615 18108 25136 18136
rect 23615 18105 23627 18108
rect 23569 18099 23627 18105
rect 25130 18096 25136 18108
rect 25188 18096 25194 18148
rect 25222 18096 25228 18148
rect 25280 18136 25286 18148
rect 26988 18136 27016 18167
rect 27706 18164 27712 18216
rect 27764 18204 27770 18216
rect 30098 18204 30104 18216
rect 27764 18176 28994 18204
rect 30059 18176 30104 18204
rect 27764 18164 27770 18176
rect 28966 18136 28994 18176
rect 30098 18164 30104 18176
rect 30156 18164 30162 18216
rect 31662 18164 31668 18216
rect 31720 18204 31726 18216
rect 34241 18207 34299 18213
rect 34241 18204 34253 18207
rect 31720 18176 34253 18204
rect 31720 18164 31726 18176
rect 34241 18173 34253 18176
rect 34287 18173 34299 18207
rect 34514 18204 34520 18216
rect 34475 18176 34520 18204
rect 34241 18167 34299 18173
rect 34514 18164 34520 18176
rect 34572 18164 34578 18216
rect 34606 18164 34612 18216
rect 34664 18204 34670 18216
rect 37292 18204 37320 18235
rect 34664 18176 37320 18204
rect 34664 18164 34670 18176
rect 32398 18136 32404 18148
rect 25280 18108 26004 18136
rect 26988 18108 28120 18136
rect 28966 18108 32404 18136
rect 25280 18096 25286 18108
rect 21284 18040 23520 18068
rect 23842 18028 23848 18080
rect 23900 18068 23906 18080
rect 24121 18071 24179 18077
rect 24121 18068 24133 18071
rect 23900 18040 24133 18068
rect 23900 18028 23906 18040
rect 24121 18037 24133 18040
rect 24167 18037 24179 18071
rect 24121 18031 24179 18037
rect 24946 18028 24952 18080
rect 25004 18068 25010 18080
rect 25976 18077 26004 18108
rect 28092 18080 28120 18108
rect 32398 18096 32404 18108
rect 32456 18096 32462 18148
rect 32674 18136 32680 18148
rect 32635 18108 32680 18136
rect 32674 18096 32680 18108
rect 32732 18096 32738 18148
rect 25777 18071 25835 18077
rect 25777 18068 25789 18071
rect 25004 18040 25789 18068
rect 25004 18028 25010 18040
rect 25777 18037 25789 18040
rect 25823 18037 25835 18071
rect 25777 18031 25835 18037
rect 25961 18071 26019 18077
rect 25961 18037 25973 18071
rect 26007 18037 26019 18071
rect 25961 18031 26019 18037
rect 26050 18028 26056 18080
rect 26108 18068 26114 18080
rect 27157 18071 27215 18077
rect 27157 18068 27169 18071
rect 26108 18040 27169 18068
rect 26108 18028 26114 18040
rect 27157 18037 27169 18040
rect 27203 18037 27215 18071
rect 27157 18031 27215 18037
rect 28074 18028 28080 18080
rect 28132 18068 28138 18080
rect 28353 18071 28411 18077
rect 28353 18068 28365 18071
rect 28132 18040 28365 18068
rect 28132 18028 28138 18040
rect 28353 18037 28365 18040
rect 28399 18068 28411 18071
rect 28442 18068 28448 18080
rect 28399 18040 28448 18068
rect 28399 18037 28411 18040
rect 28353 18031 28411 18037
rect 28442 18028 28448 18040
rect 28500 18028 28506 18080
rect 31110 18028 31116 18080
rect 31168 18068 31174 18080
rect 31297 18071 31355 18077
rect 31297 18068 31309 18071
rect 31168 18040 31309 18068
rect 31168 18028 31174 18040
rect 31297 18037 31309 18040
rect 31343 18037 31355 18071
rect 31297 18031 31355 18037
rect 32950 18028 32956 18080
rect 33008 18068 33014 18080
rect 35989 18071 36047 18077
rect 35989 18068 36001 18071
rect 33008 18040 36001 18068
rect 33008 18028 33014 18040
rect 35989 18037 36001 18040
rect 36035 18068 36047 18071
rect 36262 18068 36268 18080
rect 36035 18040 36268 18068
rect 36035 18037 36047 18040
rect 35989 18031 36047 18037
rect 36262 18028 36268 18040
rect 36320 18028 36326 18080
rect 36630 18068 36636 18080
rect 36591 18040 36636 18068
rect 36630 18028 36636 18040
rect 36688 18028 36694 18080
rect 37918 18028 37924 18080
rect 37976 18068 37982 18080
rect 38013 18071 38071 18077
rect 38013 18068 38025 18071
rect 37976 18040 38025 18068
rect 37976 18028 37982 18040
rect 38013 18037 38025 18040
rect 38059 18037 38071 18071
rect 38013 18031 38071 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 9324 17836 11192 17864
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1670 17728 1676 17740
rect 1443 17700 1676 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 9324 17669 9352 17836
rect 11164 17796 11192 17836
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 14093 17867 14151 17873
rect 14093 17864 14105 17867
rect 11296 17836 14105 17864
rect 11296 17824 11302 17836
rect 14093 17833 14105 17836
rect 14139 17833 14151 17867
rect 14093 17827 14151 17833
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 16117 17867 16175 17873
rect 16117 17864 16129 17867
rect 15896 17836 16129 17864
rect 15896 17824 15902 17836
rect 16117 17833 16129 17836
rect 16163 17833 16175 17867
rect 18598 17864 18604 17876
rect 18559 17836 18604 17864
rect 16117 17827 16175 17833
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 19242 17864 19248 17876
rect 19203 17836 19248 17864
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 19392 17836 19625 17864
rect 19392 17824 19398 17836
rect 19613 17833 19625 17836
rect 19659 17833 19671 17867
rect 19613 17827 19671 17833
rect 23201 17867 23259 17873
rect 23201 17833 23213 17867
rect 23247 17864 23259 17867
rect 23474 17864 23480 17876
rect 23247 17836 23480 17864
rect 23247 17833 23259 17836
rect 23201 17827 23259 17833
rect 23474 17824 23480 17836
rect 23532 17824 23538 17876
rect 23750 17824 23756 17876
rect 23808 17864 23814 17876
rect 24397 17867 24455 17873
rect 24397 17864 24409 17867
rect 23808 17836 24409 17864
rect 23808 17824 23814 17836
rect 24397 17833 24409 17836
rect 24443 17833 24455 17867
rect 24397 17827 24455 17833
rect 25869 17867 25927 17873
rect 25869 17833 25881 17867
rect 25915 17864 25927 17867
rect 26050 17864 26056 17876
rect 25915 17836 26056 17864
rect 25915 17833 25927 17836
rect 25869 17827 25927 17833
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 26326 17864 26332 17876
rect 26287 17836 26332 17864
rect 26326 17824 26332 17836
rect 26384 17824 26390 17876
rect 29914 17824 29920 17876
rect 29972 17864 29978 17876
rect 30101 17867 30159 17873
rect 30101 17864 30113 17867
rect 29972 17836 30113 17864
rect 29972 17824 29978 17836
rect 30101 17833 30113 17836
rect 30147 17864 30159 17867
rect 32493 17867 32551 17873
rect 30147 17836 32444 17864
rect 30147 17833 30159 17836
rect 30101 17827 30159 17833
rect 13081 17799 13139 17805
rect 13081 17796 13093 17799
rect 11164 17768 13093 17796
rect 13081 17765 13093 17768
rect 13127 17765 13139 17799
rect 13081 17759 13139 17765
rect 21821 17799 21879 17805
rect 21821 17765 21833 17799
rect 21867 17796 21879 17799
rect 24854 17796 24860 17808
rect 21867 17768 24860 17796
rect 21867 17765 21879 17768
rect 21821 17759 21879 17765
rect 24854 17756 24860 17768
rect 24912 17756 24918 17808
rect 25130 17756 25136 17808
rect 25188 17796 25194 17808
rect 25317 17799 25375 17805
rect 25317 17796 25329 17799
rect 25188 17768 25329 17796
rect 25188 17756 25194 17768
rect 25317 17765 25329 17768
rect 25363 17796 25375 17799
rect 26234 17796 26240 17808
rect 25363 17768 26240 17796
rect 25363 17765 25375 17768
rect 25317 17759 25375 17765
rect 26234 17756 26240 17768
rect 26292 17796 26298 17808
rect 30650 17796 30656 17808
rect 26292 17768 26556 17796
rect 26292 17756 26298 17768
rect 9585 17731 9643 17737
rect 9585 17697 9597 17731
rect 9631 17728 9643 17731
rect 9674 17728 9680 17740
rect 9631 17700 9680 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 10226 17688 10232 17740
rect 10284 17728 10290 17740
rect 10505 17731 10563 17737
rect 10505 17728 10517 17731
rect 10284 17700 10517 17728
rect 10284 17688 10290 17700
rect 10505 17697 10517 17700
rect 10551 17697 10563 17731
rect 14734 17728 14740 17740
rect 14695 17700 14740 17728
rect 10505 17691 10563 17697
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 17129 17731 17187 17737
rect 17129 17728 17141 17731
rect 16724 17700 17141 17728
rect 16724 17688 16730 17700
rect 17129 17697 17141 17700
rect 17175 17697 17187 17731
rect 18414 17728 18420 17740
rect 18375 17700 18420 17728
rect 17129 17691 17187 17697
rect 18414 17688 18420 17700
rect 18472 17688 18478 17740
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17728 19763 17731
rect 20346 17728 20352 17740
rect 19751 17700 20352 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 20346 17688 20352 17700
rect 20404 17688 20410 17740
rect 22370 17728 22376 17740
rect 22066 17700 22376 17728
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17660 8447 17663
rect 9309 17663 9367 17669
rect 8435 17632 8984 17660
rect 8435 17629 8447 17632
rect 8389 17623 8447 17629
rect 1581 17595 1639 17601
rect 1581 17561 1593 17595
rect 1627 17592 1639 17595
rect 1946 17592 1952 17604
rect 1627 17564 1952 17592
rect 1627 17561 1639 17564
rect 1581 17555 1639 17561
rect 1946 17552 1952 17564
rect 2004 17552 2010 17604
rect 8018 17484 8024 17536
rect 8076 17524 8082 17536
rect 8956 17533 8984 17632
rect 9309 17629 9321 17663
rect 9355 17629 9367 17663
rect 9309 17623 9367 17629
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10597 17663 10655 17669
rect 10597 17629 10609 17663
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 9401 17595 9459 17601
rect 9401 17561 9413 17595
rect 9447 17592 9459 17595
rect 9950 17592 9956 17604
rect 9447 17564 9956 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 9950 17552 9956 17564
rect 10008 17552 10014 17604
rect 8205 17527 8263 17533
rect 8205 17524 8217 17527
rect 8076 17496 8217 17524
rect 8076 17484 8082 17496
rect 8205 17493 8217 17496
rect 8251 17493 8263 17527
rect 8205 17487 8263 17493
rect 8941 17527 8999 17533
rect 8941 17493 8953 17527
rect 8987 17493 8999 17527
rect 8941 17487 8999 17493
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 10229 17527 10287 17533
rect 10229 17524 10241 17527
rect 9824 17496 10241 17524
rect 9824 17484 9830 17496
rect 10229 17493 10241 17496
rect 10275 17493 10287 17527
rect 10428 17524 10456 17623
rect 10612 17592 10640 17623
rect 10686 17620 10692 17672
rect 10744 17660 10750 17672
rect 11238 17660 11244 17672
rect 10744 17632 10789 17660
rect 11199 17632 11244 17660
rect 10744 17620 10750 17632
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11514 17660 11520 17672
rect 11427 17632 11520 17660
rect 11514 17620 11520 17632
rect 11572 17660 11578 17672
rect 12158 17660 12164 17672
rect 11572 17632 12164 17660
rect 11572 17620 11578 17632
rect 12158 17620 12164 17632
rect 12216 17660 12222 17672
rect 12897 17663 12955 17669
rect 12897 17660 12909 17663
rect 12216 17632 12909 17660
rect 12216 17620 12222 17632
rect 12897 17629 12909 17632
rect 12943 17660 12955 17663
rect 12986 17660 12992 17672
rect 12943 17632 12992 17660
rect 12943 17629 12955 17632
rect 12897 17623 12955 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13412 17632 14105 17660
rect 13412 17620 13418 17632
rect 14093 17629 14105 17632
rect 14139 17660 14151 17663
rect 14277 17663 14335 17669
rect 14139 17632 14228 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 11606 17592 11612 17604
rect 10612 17564 11612 17592
rect 11606 17552 11612 17564
rect 11664 17592 11670 17604
rect 12529 17595 12587 17601
rect 12529 17592 12541 17595
rect 11664 17564 12541 17592
rect 11664 17552 11670 17564
rect 12529 17561 12541 17564
rect 12575 17561 12587 17595
rect 12529 17555 12587 17561
rect 12805 17595 12863 17601
rect 12805 17561 12817 17595
rect 12851 17592 12863 17595
rect 13906 17592 13912 17604
rect 12851 17564 13912 17592
rect 12851 17561 12863 17564
rect 12805 17555 12863 17561
rect 13906 17552 13912 17564
rect 13964 17552 13970 17604
rect 11514 17524 11520 17536
rect 10428 17496 11520 17524
rect 10229 17487 10287 17493
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 12713 17527 12771 17533
rect 12713 17524 12725 17527
rect 11848 17496 12725 17524
rect 11848 17484 11854 17496
rect 12713 17493 12725 17496
rect 12759 17493 12771 17527
rect 14200 17524 14228 17632
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14550 17660 14556 17672
rect 14323 17632 14556 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 17218 17660 17224 17672
rect 16632 17632 17224 17660
rect 16632 17620 16638 17632
rect 17218 17620 17224 17632
rect 17276 17660 17282 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17276 17632 17417 17660
rect 17276 17620 17282 17632
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 18690 17660 18696 17672
rect 18651 17632 18696 17660
rect 17405 17623 17463 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 18966 17620 18972 17672
rect 19024 17660 19030 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 19024 17632 19441 17660
rect 19024 17620 19030 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 20625 17663 20683 17669
rect 20625 17629 20637 17663
rect 20671 17660 20683 17663
rect 21269 17663 21327 17669
rect 21269 17660 21281 17663
rect 20671 17632 21281 17660
rect 20671 17629 20683 17632
rect 20625 17623 20683 17629
rect 21269 17629 21281 17632
rect 21315 17660 21327 17663
rect 21729 17663 21787 17669
rect 21729 17660 21741 17663
rect 21315 17632 21741 17660
rect 21315 17629 21327 17632
rect 21269 17623 21327 17629
rect 21729 17629 21741 17632
rect 21775 17660 21787 17663
rect 22066 17660 22094 17700
rect 22370 17688 22376 17700
rect 22428 17728 22434 17740
rect 26528 17737 26556 17768
rect 28460 17768 30656 17796
rect 26513 17731 26571 17737
rect 22428 17700 23888 17728
rect 22428 17688 22434 17700
rect 23860 17672 23888 17700
rect 25516 17700 25912 17728
rect 21775 17632 22094 17660
rect 22557 17663 22615 17669
rect 21775 17629 21787 17632
rect 21729 17623 21787 17629
rect 22557 17629 22569 17663
rect 22603 17660 22615 17663
rect 22646 17660 22652 17672
rect 22603 17632 22652 17660
rect 22603 17629 22615 17632
rect 22557 17623 22615 17629
rect 22646 17620 22652 17632
rect 22704 17620 22710 17672
rect 23014 17660 23020 17672
rect 22975 17632 23020 17660
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 23201 17663 23259 17669
rect 23201 17629 23213 17663
rect 23247 17660 23259 17663
rect 23290 17660 23296 17672
rect 23247 17632 23296 17660
rect 23247 17629 23259 17632
rect 23201 17623 23259 17629
rect 23290 17620 23296 17632
rect 23348 17620 23354 17672
rect 23842 17660 23848 17672
rect 23803 17632 23848 17660
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24946 17660 24952 17672
rect 24627 17632 24952 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 15004 17595 15062 17601
rect 15004 17561 15016 17595
rect 15050 17592 15062 17595
rect 15194 17592 15200 17604
rect 15050 17564 15200 17592
rect 15050 17561 15062 17564
rect 15004 17555 15062 17561
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 18417 17595 18475 17601
rect 18417 17592 18429 17595
rect 16540 17564 18429 17592
rect 16540 17552 16546 17564
rect 18417 17561 18429 17564
rect 18463 17561 18475 17595
rect 18417 17555 18475 17561
rect 22465 17595 22523 17601
rect 22465 17561 22477 17595
rect 22511 17592 22523 17595
rect 23566 17592 23572 17604
rect 22511 17564 23572 17592
rect 22511 17561 22523 17564
rect 22465 17555 22523 17561
rect 23566 17552 23572 17564
rect 23624 17552 23630 17604
rect 15838 17524 15844 17536
rect 14200 17496 15844 17524
rect 12713 17487 12771 17493
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 20533 17527 20591 17533
rect 20533 17493 20545 17527
rect 20579 17524 20591 17527
rect 20714 17524 20720 17536
rect 20579 17496 20720 17524
rect 20579 17493 20591 17496
rect 20533 17487 20591 17493
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21174 17524 21180 17536
rect 21135 17496 21180 17524
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 23753 17527 23811 17533
rect 23753 17493 23765 17527
rect 23799 17524 23811 17527
rect 23842 17524 23848 17536
rect 23799 17496 23848 17524
rect 23799 17493 23811 17496
rect 23753 17487 23811 17493
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 25516 17533 25544 17700
rect 25884 17660 25912 17700
rect 26513 17697 26525 17731
rect 26559 17697 26571 17731
rect 26513 17691 26571 17697
rect 27614 17688 27620 17740
rect 27672 17728 27678 17740
rect 27672 17700 28212 17728
rect 27672 17688 27678 17700
rect 26605 17663 26663 17669
rect 26605 17660 26617 17663
rect 25884 17632 26617 17660
rect 26605 17629 26617 17632
rect 26651 17629 26663 17663
rect 26605 17623 26663 17629
rect 26878 17620 26884 17672
rect 26936 17660 26942 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26936 17632 26985 17660
rect 26936 17620 26942 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 27522 17620 27528 17672
rect 27580 17660 27586 17672
rect 28184 17669 28212 17700
rect 28460 17669 28488 17768
rect 30650 17756 30656 17768
rect 30708 17756 30714 17808
rect 32416 17796 32444 17836
rect 32493 17833 32505 17867
rect 32539 17864 32551 17867
rect 32858 17864 32864 17876
rect 32539 17836 32864 17864
rect 32539 17833 32551 17836
rect 32493 17827 32551 17833
rect 32858 17824 32864 17836
rect 32916 17864 32922 17876
rect 33042 17864 33048 17876
rect 32916 17836 33048 17864
rect 32916 17824 32922 17836
rect 33042 17824 33048 17836
rect 33100 17824 33106 17876
rect 34514 17824 34520 17876
rect 34572 17864 34578 17876
rect 34701 17867 34759 17873
rect 34701 17864 34713 17867
rect 34572 17836 34713 17864
rect 34572 17824 34578 17836
rect 34701 17833 34713 17836
rect 34747 17833 34759 17867
rect 34701 17827 34759 17833
rect 35342 17824 35348 17876
rect 35400 17864 35406 17876
rect 35529 17867 35587 17873
rect 35529 17864 35541 17867
rect 35400 17836 35541 17864
rect 35400 17824 35406 17836
rect 35529 17833 35541 17836
rect 35575 17833 35587 17867
rect 35529 17827 35587 17833
rect 32677 17799 32735 17805
rect 32416 17768 32628 17796
rect 28718 17688 28724 17740
rect 28776 17728 28782 17740
rect 32600 17728 32628 17768
rect 32677 17765 32689 17799
rect 32723 17796 32735 17799
rect 32766 17796 32772 17808
rect 32723 17768 32772 17796
rect 32723 17765 32735 17768
rect 32677 17759 32735 17765
rect 32766 17756 32772 17768
rect 32824 17796 32830 17808
rect 33229 17799 33287 17805
rect 33229 17796 33241 17799
rect 32824 17768 33241 17796
rect 32824 17756 32830 17768
rect 33229 17765 33241 17768
rect 33275 17765 33287 17799
rect 33229 17759 33287 17765
rect 33870 17756 33876 17808
rect 33928 17796 33934 17808
rect 35250 17796 35256 17808
rect 33928 17768 35256 17796
rect 33928 17756 33934 17768
rect 35250 17756 35256 17768
rect 35308 17756 35314 17808
rect 35434 17756 35440 17808
rect 35492 17796 35498 17808
rect 35621 17799 35679 17805
rect 35621 17796 35633 17799
rect 35492 17768 35633 17796
rect 35492 17756 35498 17768
rect 35621 17765 35633 17768
rect 35667 17765 35679 17799
rect 37458 17796 37464 17808
rect 35621 17759 35679 17765
rect 35728 17768 37464 17796
rect 35728 17728 35756 17768
rect 37458 17756 37464 17768
rect 37516 17756 37522 17808
rect 38010 17756 38016 17808
rect 38068 17756 38074 17808
rect 37090 17728 37096 17740
rect 28776 17700 31248 17728
rect 32600 17700 35756 17728
rect 37051 17700 37096 17728
rect 28776 17688 28782 17700
rect 27893 17663 27951 17669
rect 27893 17660 27905 17663
rect 27580 17632 27905 17660
rect 27580 17620 27586 17632
rect 27893 17629 27905 17632
rect 27939 17629 27951 17663
rect 27893 17623 27951 17629
rect 28169 17663 28227 17669
rect 28169 17629 28181 17663
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 28445 17663 28503 17669
rect 28445 17629 28457 17663
rect 28491 17629 28503 17663
rect 28445 17623 28503 17629
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17660 28687 17663
rect 29822 17660 29828 17672
rect 28675 17632 29828 17660
rect 28675 17629 28687 17632
rect 28629 17623 28687 17629
rect 29822 17620 29828 17632
rect 29880 17620 29886 17672
rect 30098 17620 30104 17672
rect 30156 17660 30162 17672
rect 31113 17663 31171 17669
rect 31113 17660 31125 17663
rect 30156 17632 31125 17660
rect 30156 17620 30162 17632
rect 31113 17629 31125 17632
rect 31159 17629 31171 17663
rect 31113 17623 31171 17629
rect 25593 17595 25651 17601
rect 25593 17561 25605 17595
rect 25639 17592 25651 17595
rect 27706 17592 27712 17604
rect 25639 17564 26740 17592
rect 25639 17561 25651 17564
rect 25593 17555 25651 17561
rect 26712 17536 26740 17564
rect 26896 17564 27712 17592
rect 25501 17527 25559 17533
rect 25501 17524 25513 17527
rect 24636 17496 25513 17524
rect 24636 17484 24642 17496
rect 25501 17493 25513 17496
rect 25547 17493 25559 17527
rect 25501 17487 25559 17493
rect 25685 17527 25743 17533
rect 25685 17493 25697 17527
rect 25731 17524 25743 17527
rect 26510 17524 26516 17536
rect 25731 17496 26516 17524
rect 25731 17493 25743 17496
rect 25685 17487 25743 17493
rect 26510 17484 26516 17496
rect 26568 17484 26574 17536
rect 26694 17524 26700 17536
rect 26607 17496 26700 17524
rect 26694 17484 26700 17496
rect 26752 17484 26758 17536
rect 26896 17533 26924 17564
rect 27706 17552 27712 17564
rect 27764 17552 27770 17604
rect 28258 17552 28264 17604
rect 28316 17592 28322 17604
rect 30009 17595 30067 17601
rect 30009 17592 30021 17595
rect 28316 17564 30021 17592
rect 28316 17552 28322 17564
rect 30009 17561 30021 17564
rect 30055 17561 30067 17595
rect 31220 17592 31248 17700
rect 33137 17663 33195 17669
rect 33137 17629 33149 17663
rect 33183 17660 33195 17663
rect 33226 17660 33232 17672
rect 33183 17632 33232 17660
rect 33183 17629 33195 17632
rect 33137 17623 33195 17629
rect 33226 17620 33232 17632
rect 33284 17620 33290 17672
rect 33428 17669 33456 17700
rect 37090 17688 37096 17700
rect 37148 17688 37154 17740
rect 37918 17728 37924 17740
rect 37879 17700 37924 17728
rect 37918 17688 37924 17700
rect 37976 17688 37982 17740
rect 38028 17728 38056 17756
rect 38105 17731 38163 17737
rect 38105 17728 38117 17731
rect 38028 17700 38117 17728
rect 38105 17697 38117 17700
rect 38151 17697 38163 17731
rect 38105 17691 38163 17697
rect 33413 17663 33471 17669
rect 33413 17629 33425 17663
rect 33459 17629 33471 17663
rect 33413 17623 33471 17629
rect 33686 17620 33692 17672
rect 33744 17660 33750 17672
rect 34977 17663 35035 17669
rect 34977 17660 34989 17663
rect 33744 17632 34989 17660
rect 33744 17620 33750 17632
rect 34977 17629 34989 17632
rect 35023 17629 35035 17663
rect 34977 17623 35035 17629
rect 35250 17620 35256 17672
rect 35308 17660 35314 17672
rect 35437 17663 35495 17669
rect 35437 17660 35449 17663
rect 35308 17632 35449 17660
rect 35308 17620 35314 17632
rect 35437 17629 35449 17632
rect 35483 17660 35495 17663
rect 35526 17660 35532 17672
rect 35483 17632 35532 17660
rect 35483 17629 35495 17632
rect 35437 17623 35495 17629
rect 35526 17620 35532 17632
rect 35584 17620 35590 17672
rect 35713 17663 35771 17669
rect 35713 17629 35725 17663
rect 35759 17660 35771 17663
rect 35802 17660 35808 17672
rect 35759 17632 35808 17660
rect 35759 17629 35771 17632
rect 35713 17623 35771 17629
rect 35802 17620 35808 17632
rect 35860 17620 35866 17672
rect 32309 17595 32367 17601
rect 31220 17564 31754 17592
rect 30009 17555 30067 17561
rect 26881 17527 26939 17533
rect 26881 17493 26893 17527
rect 26927 17493 26939 17527
rect 26881 17487 26939 17493
rect 27154 17484 27160 17536
rect 27212 17524 27218 17536
rect 27985 17527 28043 17533
rect 27985 17524 27997 17527
rect 27212 17496 27997 17524
rect 27212 17484 27218 17496
rect 27985 17493 27997 17496
rect 28031 17493 28043 17527
rect 27985 17487 28043 17493
rect 30742 17484 30748 17536
rect 30800 17524 30806 17536
rect 31205 17527 31263 17533
rect 31205 17524 31217 17527
rect 30800 17496 31217 17524
rect 30800 17484 30806 17496
rect 31205 17493 31217 17496
rect 31251 17524 31263 17527
rect 31386 17524 31392 17536
rect 31251 17496 31392 17524
rect 31251 17493 31263 17496
rect 31205 17487 31263 17493
rect 31386 17484 31392 17496
rect 31444 17484 31450 17536
rect 31726 17524 31754 17564
rect 32309 17561 32321 17595
rect 32355 17592 32367 17595
rect 32950 17592 32956 17604
rect 32355 17564 32956 17592
rect 32355 17561 32367 17564
rect 32309 17555 32367 17561
rect 32950 17552 32956 17564
rect 33008 17552 33014 17604
rect 33597 17595 33655 17601
rect 33597 17561 33609 17595
rect 33643 17592 33655 17595
rect 34701 17595 34759 17601
rect 34701 17592 34713 17595
rect 33643 17564 34713 17592
rect 33643 17561 33655 17564
rect 33597 17555 33655 17561
rect 34701 17561 34713 17564
rect 34747 17561 34759 17595
rect 34701 17555 34759 17561
rect 32398 17524 32404 17536
rect 31726 17496 32404 17524
rect 32398 17484 32404 17496
rect 32456 17484 32462 17536
rect 32490 17484 32496 17536
rect 32548 17533 32554 17536
rect 32548 17527 32567 17533
rect 32555 17493 32567 17527
rect 34882 17524 34888 17536
rect 34843 17496 34888 17524
rect 32548 17487 32567 17493
rect 32548 17484 32554 17487
rect 34882 17484 34888 17496
rect 34940 17484 34946 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9674 17320 9680 17332
rect 9171 17292 9680 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 10560 17292 10701 17320
rect 10560 17280 10566 17292
rect 10689 17289 10701 17292
rect 10735 17289 10747 17323
rect 10689 17283 10747 17289
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 14550 17320 14556 17332
rect 10836 17292 10881 17320
rect 14511 17292 14556 17320
rect 10836 17280 10842 17292
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 15194 17320 15200 17332
rect 15155 17292 15200 17320
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 16666 17320 16672 17332
rect 16627 17292 16672 17320
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 18693 17323 18751 17329
rect 18693 17289 18705 17323
rect 18739 17320 18751 17323
rect 18966 17320 18972 17332
rect 18739 17292 18972 17320
rect 18739 17289 18751 17292
rect 18693 17283 18751 17289
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 22465 17323 22523 17329
rect 22465 17289 22477 17323
rect 22511 17320 22523 17323
rect 22554 17320 22560 17332
rect 22511 17292 22560 17320
rect 22511 17289 22523 17292
rect 22465 17283 22523 17289
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 27154 17320 27160 17332
rect 24728 17292 27160 17320
rect 24728 17280 24734 17292
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 27522 17320 27528 17332
rect 27483 17292 27528 17320
rect 27522 17280 27528 17292
rect 27580 17280 27586 17332
rect 27614 17280 27620 17332
rect 27672 17320 27678 17332
rect 32030 17320 32036 17332
rect 27672 17292 32036 17320
rect 27672 17280 27678 17292
rect 32030 17280 32036 17292
rect 32088 17280 32094 17332
rect 32858 17329 32864 17332
rect 32845 17323 32864 17329
rect 32845 17289 32857 17323
rect 32845 17283 32864 17289
rect 32858 17280 32864 17283
rect 32916 17280 32922 17332
rect 33134 17280 33140 17332
rect 33192 17320 33198 17332
rect 33705 17323 33763 17329
rect 33705 17320 33717 17323
rect 33192 17292 33717 17320
rect 33192 17280 33198 17292
rect 33705 17289 33717 17292
rect 33751 17289 33763 17323
rect 33705 17283 33763 17289
rect 33873 17323 33931 17329
rect 33873 17289 33885 17323
rect 33919 17320 33931 17323
rect 34606 17320 34612 17332
rect 33919 17292 34612 17320
rect 33919 17289 33931 17292
rect 33873 17283 33931 17289
rect 34606 17280 34612 17292
rect 34664 17280 34670 17332
rect 34882 17280 34888 17332
rect 34940 17320 34946 17332
rect 37369 17323 37427 17329
rect 37369 17320 37381 17323
rect 34940 17292 37381 17320
rect 34940 17280 34946 17292
rect 37369 17289 37381 17292
rect 37415 17289 37427 17323
rect 37369 17283 37427 17289
rect 8662 17252 8668 17264
rect 7760 17224 8668 17252
rect 2038 17184 2044 17196
rect 1999 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 7760 17193 7788 17224
rect 8662 17212 8668 17224
rect 8720 17212 8726 17264
rect 13633 17255 13691 17261
rect 13633 17221 13645 17255
rect 13679 17252 13691 17255
rect 13998 17252 14004 17264
rect 13679 17224 14004 17252
rect 13679 17221 13691 17224
rect 13633 17215 13691 17221
rect 13998 17212 14004 17224
rect 14056 17252 14062 17264
rect 14056 17224 14780 17252
rect 14056 17212 14062 17224
rect 8018 17193 8024 17196
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17153 7803 17187
rect 8012 17184 8024 17193
rect 7979 17156 8024 17184
rect 7745 17147 7803 17153
rect 8012 17147 8024 17156
rect 8018 17144 8024 17147
rect 8076 17144 8082 17196
rect 9766 17184 9772 17196
rect 9727 17156 9772 17184
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 11238 17184 11244 17196
rect 10919 17156 11244 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11664 17156 11805 17184
rect 11664 17144 11670 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 11793 17147 11851 17153
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 13078 17144 13084 17196
rect 13136 17184 13142 17196
rect 14752 17193 14780 17224
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 16025 17255 16083 17261
rect 15344 17224 15976 17252
rect 15344 17212 15350 17224
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13136 17156 13921 17184
rect 13136 17144 13142 17156
rect 13909 17153 13921 17156
rect 13955 17184 13967 17187
rect 14553 17187 14611 17193
rect 14553 17184 14565 17187
rect 13955 17156 14565 17184
rect 13955 17153 13967 17156
rect 13909 17147 13967 17153
rect 14553 17153 14565 17156
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17153 14795 17187
rect 15378 17184 15384 17196
rect 15339 17156 15384 17184
rect 14737 17147 14795 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 15948 17193 15976 17224
rect 16025 17221 16037 17255
rect 16071 17252 16083 17255
rect 18138 17252 18144 17264
rect 16071 17224 18144 17252
rect 16071 17221 16083 17224
rect 16025 17215 16083 17221
rect 18138 17212 18144 17224
rect 18196 17212 18202 17264
rect 18414 17212 18420 17264
rect 18472 17252 18478 17264
rect 21174 17252 21180 17264
rect 18472 17224 18736 17252
rect 21022 17224 21180 17252
rect 18472 17212 18478 17224
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17184 16175 17187
rect 16298 17184 16304 17196
rect 16163 17156 16304 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17782 17187 17840 17193
rect 17782 17184 17794 17187
rect 17000 17156 17794 17184
rect 17000 17144 17006 17156
rect 17782 17153 17794 17156
rect 17828 17153 17840 17187
rect 17782 17147 17840 17153
rect 17954 17144 17960 17196
rect 18012 17184 18018 17196
rect 18049 17187 18107 17193
rect 18049 17184 18061 17187
rect 18012 17156 18061 17184
rect 18012 17144 18018 17156
rect 18049 17153 18061 17156
rect 18095 17153 18107 17187
rect 18506 17184 18512 17196
rect 18467 17156 18512 17184
rect 18049 17147 18107 17153
rect 9950 17116 9956 17128
rect 9911 17088 9956 17116
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17116 10563 17119
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 10551 17088 11529 17116
rect 10551 17085 10563 17088
rect 10505 17079 10563 17085
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 13173 17119 13231 17125
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13446 17116 13452 17128
rect 13219 17088 13452 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 10781 17051 10839 17057
rect 10781 17017 10793 17051
rect 10827 17048 10839 17051
rect 10962 17048 10968 17060
rect 10827 17020 10968 17048
rect 10827 17017 10839 17020
rect 10781 17011 10839 17017
rect 10962 17008 10968 17020
rect 11020 17008 11026 17060
rect 11532 17048 11560 17079
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17085 13783 17119
rect 18064 17116 18092 17147
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18708 17193 18736 17224
rect 21174 17212 21180 17224
rect 21232 17212 21238 17264
rect 23842 17212 23848 17264
rect 23900 17212 23906 17264
rect 27065 17255 27123 17261
rect 27065 17221 27077 17255
rect 27111 17252 27123 17255
rect 27246 17252 27252 17264
rect 27111 17224 27252 17252
rect 27111 17221 27123 17224
rect 27065 17215 27123 17221
rect 27246 17212 27252 17224
rect 27304 17212 27310 17264
rect 27430 17212 27436 17264
rect 27488 17252 27494 17264
rect 27488 17224 29946 17252
rect 27488 17212 27494 17224
rect 32674 17212 32680 17264
rect 32732 17252 32738 17264
rect 33042 17252 33048 17264
rect 32732 17224 33048 17252
rect 32732 17212 32738 17224
rect 33042 17212 33048 17224
rect 33100 17212 33106 17264
rect 33505 17255 33563 17261
rect 33505 17221 33517 17255
rect 33551 17252 33563 17255
rect 33594 17252 33600 17264
rect 33551 17224 33600 17252
rect 33551 17221 33563 17224
rect 33505 17215 33563 17221
rect 33594 17212 33600 17224
rect 33652 17212 33658 17264
rect 35069 17255 35127 17261
rect 35069 17221 35081 17255
rect 35115 17252 35127 17255
rect 38013 17255 38071 17261
rect 38013 17252 38025 17255
rect 35115 17224 38025 17252
rect 35115 17221 35127 17224
rect 35069 17215 35127 17221
rect 38013 17221 38025 17224
rect 38059 17221 38071 17255
rect 38013 17215 38071 17221
rect 18693 17187 18751 17193
rect 18693 17153 18705 17187
rect 18739 17153 18751 17187
rect 22370 17184 22376 17196
rect 22331 17156 22376 17184
rect 18693 17147 18751 17153
rect 22370 17144 22376 17156
rect 22428 17144 22434 17196
rect 24857 17187 24915 17193
rect 24857 17153 24869 17187
rect 24903 17184 24915 17187
rect 25038 17184 25044 17196
rect 24903 17156 25044 17184
rect 24903 17153 24915 17156
rect 24857 17147 24915 17153
rect 25038 17144 25044 17156
rect 25096 17144 25102 17196
rect 25498 17184 25504 17196
rect 25459 17156 25504 17184
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 25593 17187 25651 17193
rect 25593 17153 25605 17187
rect 25639 17153 25651 17187
rect 25593 17147 25651 17153
rect 19426 17116 19432 17128
rect 18064 17088 19432 17116
rect 13725 17079 13783 17085
rect 12894 17048 12900 17060
rect 11532 17020 12900 17048
rect 12894 17008 12900 17020
rect 12952 17048 12958 17060
rect 13740 17048 13768 17079
rect 19426 17076 19432 17088
rect 19484 17116 19490 17128
rect 19521 17119 19579 17125
rect 19521 17116 19533 17119
rect 19484 17088 19533 17116
rect 19484 17076 19490 17088
rect 19521 17085 19533 17088
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 19797 17119 19855 17125
rect 19797 17085 19809 17119
rect 19843 17116 19855 17119
rect 20162 17116 20168 17128
rect 19843 17088 20168 17116
rect 19843 17085 19855 17088
rect 19797 17079 19855 17085
rect 20162 17076 20168 17088
rect 20220 17076 20226 17128
rect 24581 17119 24639 17125
rect 24581 17085 24593 17119
rect 24627 17116 24639 17119
rect 25608 17116 25636 17147
rect 25682 17144 25688 17196
rect 25740 17184 25746 17196
rect 25740 17156 25785 17184
rect 25740 17144 25746 17156
rect 25866 17144 25872 17196
rect 25924 17184 25930 17196
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 25924 17156 25969 17184
rect 26988 17156 27353 17184
rect 25924 17144 25930 17156
rect 26988 17116 27016 17156
rect 27341 17153 27353 17156
rect 27387 17153 27399 17187
rect 28258 17184 28264 17196
rect 28219 17156 28264 17184
rect 27341 17147 27399 17153
rect 28258 17144 28264 17156
rect 28316 17144 28322 17196
rect 36262 17144 36268 17196
rect 36320 17184 36326 17196
rect 37277 17187 37335 17193
rect 37277 17184 37289 17187
rect 36320 17156 37289 17184
rect 36320 17144 36326 17156
rect 37277 17153 37289 17156
rect 37323 17153 37335 17187
rect 37277 17147 37335 17153
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17153 37979 17187
rect 37921 17147 37979 17153
rect 24627 17088 25360 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 12952 17020 13768 17048
rect 14093 17051 14151 17057
rect 12952 17008 12958 17020
rect 14093 17017 14105 17051
rect 14139 17048 14151 17051
rect 14826 17048 14832 17060
rect 14139 17020 14832 17048
rect 14139 17017 14151 17020
rect 14093 17011 14151 17017
rect 14826 17008 14832 17020
rect 14884 17008 14890 17060
rect 25332 17057 25360 17088
rect 25608 17088 27016 17116
rect 27249 17119 27307 17125
rect 25317 17051 25375 17057
rect 25317 17017 25329 17051
rect 25363 17017 25375 17051
rect 25317 17011 25375 17017
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 9456 16952 9597 16980
rect 9456 16940 9462 16952
rect 9585 16949 9597 16952
rect 9631 16949 9643 16983
rect 9585 16943 9643 16949
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12676 16952 12817 16980
rect 12676 16940 12682 16952
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 13722 16980 13728 16992
rect 13683 16952 13728 16980
rect 12805 16943 12863 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21269 16983 21327 16989
rect 21269 16980 21281 16983
rect 20956 16952 21281 16980
rect 20956 16940 20962 16952
rect 21269 16949 21281 16952
rect 21315 16949 21327 16983
rect 21269 16943 21327 16949
rect 23109 16983 23167 16989
rect 23109 16949 23121 16983
rect 23155 16980 23167 16983
rect 24578 16980 24584 16992
rect 23155 16952 24584 16980
rect 23155 16949 23167 16952
rect 23109 16943 23167 16949
rect 24578 16940 24584 16952
rect 24636 16980 24642 16992
rect 25608 16980 25636 17088
rect 27249 17085 27261 17119
rect 27295 17085 27307 17119
rect 27249 17079 27307 17085
rect 25866 17008 25872 17060
rect 25924 17048 25930 17060
rect 27264 17048 27292 17079
rect 27614 17076 27620 17128
rect 27672 17116 27678 17128
rect 27985 17119 28043 17125
rect 27985 17116 27997 17119
rect 27672 17088 27997 17116
rect 27672 17076 27678 17088
rect 27985 17085 27997 17088
rect 28031 17085 28043 17119
rect 31110 17116 31116 17128
rect 31071 17088 31116 17116
rect 27985 17079 28043 17085
rect 31110 17076 31116 17088
rect 31168 17076 31174 17128
rect 31389 17119 31447 17125
rect 31389 17085 31401 17119
rect 31435 17116 31447 17119
rect 31662 17116 31668 17128
rect 31435 17088 31668 17116
rect 31435 17085 31447 17088
rect 31389 17079 31447 17085
rect 31662 17076 31668 17088
rect 31720 17076 31726 17128
rect 34885 17119 34943 17125
rect 34885 17085 34897 17119
rect 34931 17116 34943 17119
rect 35710 17116 35716 17128
rect 34931 17088 35716 17116
rect 34931 17085 34943 17088
rect 34885 17079 34943 17085
rect 35710 17076 35716 17088
rect 35768 17076 35774 17128
rect 36722 17116 36728 17128
rect 36683 17088 36728 17116
rect 36722 17076 36728 17088
rect 36780 17076 36786 17128
rect 29638 17048 29644 17060
rect 25924 17020 27200 17048
rect 27264 17020 29644 17048
rect 25924 17008 25930 17020
rect 24636 16952 25636 16980
rect 24636 16940 24642 16952
rect 26694 16940 26700 16992
rect 26752 16980 26758 16992
rect 27065 16983 27123 16989
rect 27065 16980 27077 16983
rect 26752 16952 27077 16980
rect 26752 16940 26758 16952
rect 27065 16949 27077 16952
rect 27111 16949 27123 16983
rect 27172 16980 27200 17020
rect 29638 17008 29644 17020
rect 29696 17008 29702 17060
rect 32398 17008 32404 17060
rect 32456 17048 32462 17060
rect 37936 17048 37964 17147
rect 32456 17020 37964 17048
rect 32456 17008 32462 17020
rect 30742 16980 30748 16992
rect 27172 16952 30748 16980
rect 27065 16943 27123 16949
rect 30742 16940 30748 16952
rect 30800 16940 30806 16992
rect 32122 16940 32128 16992
rect 32180 16980 32186 16992
rect 32677 16983 32735 16989
rect 32677 16980 32689 16983
rect 32180 16952 32689 16980
rect 32180 16940 32186 16952
rect 32677 16949 32689 16952
rect 32723 16949 32735 16983
rect 32677 16943 32735 16949
rect 32861 16983 32919 16989
rect 32861 16949 32873 16983
rect 32907 16980 32919 16983
rect 32950 16980 32956 16992
rect 32907 16952 32956 16980
rect 32907 16949 32919 16952
rect 32861 16943 32919 16949
rect 32950 16940 32956 16952
rect 33008 16940 33014 16992
rect 33686 16980 33692 16992
rect 33647 16952 33692 16980
rect 33686 16940 33692 16952
rect 33744 16940 33750 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 10321 16779 10379 16785
rect 10321 16745 10333 16779
rect 10367 16776 10379 16779
rect 10686 16776 10692 16788
rect 10367 16748 10692 16776
rect 10367 16745 10379 16748
rect 10321 16739 10379 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 16942 16776 16948 16788
rect 16903 16748 16948 16776
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 22738 16776 22744 16788
rect 19392 16748 22744 16776
rect 19392 16736 19398 16748
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 24857 16779 24915 16785
rect 24857 16745 24869 16779
rect 24903 16776 24915 16779
rect 25682 16776 25688 16788
rect 24903 16748 25688 16776
rect 24903 16745 24915 16748
rect 24857 16739 24915 16745
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 26881 16779 26939 16785
rect 26881 16745 26893 16779
rect 26927 16776 26939 16779
rect 27798 16776 27804 16788
rect 26927 16748 27804 16776
rect 26927 16745 26939 16748
rect 26881 16739 26939 16745
rect 27798 16736 27804 16748
rect 27856 16736 27862 16788
rect 28000 16748 28994 16776
rect 11974 16708 11980 16720
rect 11624 16680 11980 16708
rect 8662 16600 8668 16652
rect 8720 16640 8726 16652
rect 11624 16649 11652 16680
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 13078 16708 13084 16720
rect 12912 16680 13084 16708
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8720 16612 8953 16640
rect 8720 16600 8726 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 11609 16643 11667 16649
rect 11609 16609 11621 16643
rect 11655 16609 11667 16643
rect 11609 16603 11667 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12912 16649 12940 16680
rect 13078 16668 13084 16680
rect 13136 16668 13142 16720
rect 15746 16668 15752 16720
rect 15804 16708 15810 16720
rect 22370 16708 22376 16720
rect 15804 16680 17448 16708
rect 22331 16680 22376 16708
rect 15804 16668 15810 16680
rect 12897 16643 12955 16649
rect 11756 16612 11801 16640
rect 11756 16600 11762 16612
rect 12897 16609 12909 16643
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 13262 16640 13268 16652
rect 13035 16612 13268 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 15933 16643 15991 16649
rect 15933 16640 15945 16643
rect 14200 16612 15945 16640
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16572 11575 16575
rect 12618 16572 12624 16584
rect 11563 16544 12624 16572
rect 11563 16541 11575 16544
rect 11517 16535 11575 16541
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16572 13139 16575
rect 14200 16572 14228 16612
rect 14660 16581 14688 16612
rect 15933 16609 15945 16612
rect 15979 16609 15991 16643
rect 17034 16640 17040 16652
rect 15933 16603 15991 16609
rect 16040 16612 17040 16640
rect 13127 16544 14228 16572
rect 14277 16575 14335 16581
rect 13127 16541 13139 16544
rect 13081 16535 13139 16541
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16541 14703 16575
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 14645 16535 14703 16541
rect 9214 16513 9220 16516
rect 9208 16467 9220 16513
rect 9272 16504 9278 16516
rect 9272 16476 9308 16504
rect 9214 16464 9220 16467
rect 9272 16464 9278 16476
rect 11974 16464 11980 16516
rect 12032 16504 12038 16516
rect 14292 16504 14320 16535
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 16040 16581 16068 16612
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 17420 16640 17448 16680
rect 22370 16668 22376 16680
rect 22428 16708 22434 16720
rect 23198 16708 23204 16720
rect 22428 16680 23204 16708
rect 22428 16668 22434 16680
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 23845 16711 23903 16717
rect 23845 16677 23857 16711
rect 23891 16708 23903 16711
rect 27522 16708 27528 16720
rect 23891 16680 27528 16708
rect 23891 16677 23903 16680
rect 23845 16671 23903 16677
rect 27522 16668 27528 16680
rect 27580 16668 27586 16720
rect 27706 16668 27712 16720
rect 27764 16708 27770 16720
rect 27890 16708 27896 16720
rect 27764 16680 27896 16708
rect 27764 16668 27770 16680
rect 27890 16668 27896 16680
rect 27948 16668 27954 16720
rect 17420 16612 18092 16640
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16482 16572 16488 16584
rect 16443 16544 16488 16572
rect 16025 16535 16083 16541
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 16574 16532 16580 16584
rect 16632 16572 16638 16584
rect 16758 16572 16764 16584
rect 16632 16544 16677 16572
rect 16719 16544 16764 16572
rect 16632 16532 16638 16544
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17420 16581 17448 16612
rect 18064 16581 18092 16612
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19484 16612 19993 16640
rect 19484 16600 19490 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 20254 16640 20260 16652
rect 20215 16612 20260 16640
rect 19981 16603 20039 16609
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22462 16640 22468 16652
rect 22152 16612 22468 16640
rect 22152 16600 22158 16612
rect 22462 16600 22468 16612
rect 22520 16640 22526 16652
rect 22557 16643 22615 16649
rect 22557 16640 22569 16643
rect 22520 16612 22569 16640
rect 22520 16600 22526 16612
rect 22557 16609 22569 16612
rect 22603 16609 22615 16643
rect 25501 16643 25559 16649
rect 25501 16640 25513 16643
rect 22557 16603 22615 16609
rect 24872 16612 25513 16640
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16541 19579 16575
rect 19521 16535 19579 16541
rect 12032 16476 14320 16504
rect 14369 16507 14427 16513
rect 12032 16464 12038 16476
rect 14369 16473 14381 16507
rect 14415 16473 14427 16507
rect 14369 16467 14427 16473
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 10836 16408 11161 16436
rect 10836 16396 10842 16408
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 11149 16399 11207 16405
rect 13170 16396 13176 16448
rect 13228 16436 13234 16448
rect 13449 16439 13507 16445
rect 13449 16436 13461 16439
rect 13228 16408 13461 16436
rect 13228 16396 13234 16408
rect 13449 16405 13461 16408
rect 13495 16405 13507 16439
rect 13449 16399 13507 16405
rect 13906 16396 13912 16448
rect 13964 16436 13970 16448
rect 14093 16439 14151 16445
rect 14093 16436 14105 16439
rect 13964 16408 14105 16436
rect 13964 16396 13970 16408
rect 14093 16405 14105 16408
rect 14139 16405 14151 16439
rect 14093 16399 14151 16405
rect 14182 16396 14188 16448
rect 14240 16436 14246 16448
rect 14384 16436 14412 16467
rect 14458 16464 14464 16516
rect 14516 16504 14522 16516
rect 19536 16504 19564 16535
rect 22186 16532 22192 16584
rect 22244 16572 22250 16584
rect 22281 16575 22339 16581
rect 22281 16572 22293 16575
rect 22244 16544 22293 16572
rect 22244 16532 22250 16544
rect 22281 16541 22293 16544
rect 22327 16541 22339 16575
rect 23198 16572 23204 16584
rect 23159 16544 23204 16572
rect 22281 16535 22339 16541
rect 23198 16532 23204 16544
rect 23256 16532 23262 16584
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23586 16575 23644 16581
rect 23586 16541 23598 16575
rect 23632 16572 23644 16575
rect 24578 16572 24584 16584
rect 23632 16544 23704 16572
rect 24539 16544 24584 16572
rect 23632 16541 23644 16544
rect 23586 16535 23644 16541
rect 20530 16504 20536 16516
rect 14516 16476 14561 16504
rect 19536 16476 20536 16504
rect 14516 16464 14522 16476
rect 20530 16464 20536 16476
rect 20588 16464 20594 16516
rect 20714 16464 20720 16516
rect 20772 16464 20778 16516
rect 22557 16507 22615 16513
rect 22557 16473 22569 16507
rect 22603 16504 22615 16507
rect 23106 16504 23112 16516
rect 22603 16476 23112 16504
rect 22603 16473 22615 16476
rect 22557 16467 22615 16473
rect 23106 16464 23112 16476
rect 23164 16504 23170 16516
rect 23400 16504 23428 16535
rect 23164 16476 23428 16504
rect 23164 16464 23170 16476
rect 14240 16408 14412 16436
rect 17497 16439 17555 16445
rect 14240 16396 14246 16408
rect 17497 16405 17509 16439
rect 17543 16436 17555 16439
rect 17954 16436 17960 16448
rect 17543 16408 17960 16436
rect 17543 16405 17555 16408
rect 17497 16399 17555 16405
rect 17954 16396 17960 16408
rect 18012 16396 18018 16448
rect 18138 16436 18144 16448
rect 18099 16408 18144 16436
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 19337 16439 19395 16445
rect 19337 16405 19349 16439
rect 19383 16436 19395 16439
rect 20070 16436 20076 16448
rect 19383 16408 20076 16436
rect 19383 16405 19395 16408
rect 19337 16399 19395 16405
rect 20070 16396 20076 16408
rect 20128 16436 20134 16448
rect 20438 16436 20444 16448
rect 20128 16408 20444 16436
rect 20128 16396 20134 16408
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 21082 16396 21088 16448
rect 21140 16436 21146 16448
rect 21729 16439 21787 16445
rect 21729 16436 21741 16439
rect 21140 16408 21741 16436
rect 21140 16396 21146 16408
rect 21729 16405 21741 16408
rect 21775 16405 21787 16439
rect 21729 16399 21787 16405
rect 22922 16396 22928 16448
rect 22980 16436 22986 16448
rect 23290 16436 23296 16448
rect 22980 16408 23296 16436
rect 22980 16396 22986 16408
rect 23290 16396 23296 16408
rect 23348 16436 23354 16448
rect 23492 16436 23520 16535
rect 23676 16504 23704 16544
rect 24578 16532 24584 16544
rect 24636 16532 24642 16584
rect 24762 16572 24768 16584
rect 24723 16544 24768 16572
rect 24762 16532 24768 16544
rect 24820 16532 24826 16584
rect 24872 16581 24900 16612
rect 25501 16609 25513 16612
rect 25547 16640 25559 16643
rect 25866 16640 25872 16652
rect 25547 16612 25872 16640
rect 25547 16609 25559 16612
rect 25501 16603 25559 16609
rect 25866 16600 25872 16612
rect 25924 16600 25930 16652
rect 26970 16600 26976 16652
rect 27028 16640 27034 16652
rect 28000 16640 28028 16748
rect 28074 16668 28080 16720
rect 28132 16708 28138 16720
rect 28966 16708 28994 16748
rect 29638 16736 29644 16788
rect 29696 16776 29702 16788
rect 29696 16748 30236 16776
rect 29696 16736 29702 16748
rect 30208 16720 30236 16748
rect 30282 16736 30288 16788
rect 30340 16776 30346 16788
rect 31205 16779 31263 16785
rect 31205 16776 31217 16779
rect 30340 16748 31217 16776
rect 30340 16736 30346 16748
rect 31205 16745 31217 16748
rect 31251 16745 31263 16779
rect 32122 16776 32128 16788
rect 32083 16748 32128 16776
rect 31205 16739 31263 16745
rect 32122 16736 32128 16748
rect 32180 16736 32186 16788
rect 33870 16776 33876 16788
rect 33831 16748 33876 16776
rect 33870 16736 33876 16748
rect 33928 16736 33934 16788
rect 34698 16776 34704 16788
rect 34659 16748 34704 16776
rect 34698 16736 34704 16748
rect 34756 16736 34762 16788
rect 35161 16779 35219 16785
rect 35161 16745 35173 16779
rect 35207 16776 35219 16779
rect 35342 16776 35348 16788
rect 35207 16748 35348 16776
rect 35207 16745 35219 16748
rect 35161 16739 35219 16745
rect 35342 16736 35348 16748
rect 35400 16736 35406 16788
rect 29362 16708 29368 16720
rect 28132 16680 28489 16708
rect 28966 16680 29368 16708
rect 28132 16668 28138 16680
rect 28461 16649 28489 16680
rect 29362 16668 29368 16680
rect 29420 16708 29426 16720
rect 29420 16680 30144 16708
rect 29420 16668 29426 16680
rect 28353 16643 28411 16649
rect 28353 16640 28365 16643
rect 27028 16612 27073 16640
rect 27422 16612 28365 16640
rect 27028 16600 27034 16612
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 25406 16532 25412 16584
rect 25464 16572 25470 16584
rect 25593 16575 25651 16581
rect 25593 16572 25605 16575
rect 25464 16544 25605 16572
rect 25464 16532 25470 16544
rect 25593 16541 25605 16544
rect 25639 16541 25651 16575
rect 25593 16535 25651 16541
rect 26142 16532 26148 16584
rect 26200 16572 26206 16584
rect 26697 16575 26755 16581
rect 26697 16572 26709 16575
rect 26200 16544 26709 16572
rect 26200 16532 26206 16544
rect 26697 16541 26709 16544
rect 26743 16541 26755 16575
rect 26697 16535 26755 16541
rect 26789 16575 26847 16581
rect 26789 16541 26801 16575
rect 26835 16572 26847 16575
rect 27422 16572 27450 16612
rect 28353 16609 28365 16612
rect 28399 16609 28411 16643
rect 28353 16603 28411 16609
rect 28445 16643 28503 16649
rect 28445 16609 28457 16643
rect 28491 16609 28503 16643
rect 28445 16603 28503 16609
rect 28626 16600 28632 16652
rect 28684 16640 28690 16652
rect 29638 16640 29644 16652
rect 28684 16612 29644 16640
rect 28684 16600 28690 16612
rect 29638 16600 29644 16612
rect 29696 16600 29702 16652
rect 27522 16572 27528 16584
rect 26835 16544 27450 16572
rect 27483 16544 27528 16572
rect 26835 16541 26847 16544
rect 26789 16535 26847 16541
rect 27522 16532 27528 16544
rect 27580 16532 27586 16584
rect 28538 16575 28596 16581
rect 28538 16566 28550 16575
rect 28461 16541 28550 16566
rect 28584 16541 28596 16575
rect 29178 16572 29184 16584
rect 28461 16538 28596 16541
rect 24486 16504 24492 16516
rect 23676 16476 24492 16504
rect 24486 16464 24492 16476
rect 24544 16464 24550 16516
rect 26160 16504 26188 16532
rect 24872 16476 26188 16504
rect 24872 16448 24900 16476
rect 27706 16464 27712 16516
rect 27764 16504 27770 16516
rect 28461 16504 28489 16538
rect 28538 16535 28596 16538
rect 28920 16544 29184 16572
rect 28920 16504 28948 16544
rect 29178 16532 29184 16544
rect 29236 16532 29242 16584
rect 30116 16581 30144 16680
rect 30190 16668 30196 16720
rect 30248 16708 30254 16720
rect 31938 16708 31944 16720
rect 30248 16680 30341 16708
rect 31899 16680 31944 16708
rect 30248 16668 30254 16680
rect 31938 16668 31944 16680
rect 31996 16668 32002 16720
rect 34057 16711 34115 16717
rect 34057 16677 34069 16711
rect 34103 16708 34115 16711
rect 37458 16708 37464 16720
rect 34103 16680 37464 16708
rect 34103 16677 34115 16680
rect 34057 16671 34115 16677
rect 37458 16668 37464 16680
rect 37516 16668 37522 16720
rect 30208 16640 30236 16668
rect 30561 16643 30619 16649
rect 30561 16640 30573 16643
rect 30208 16612 30573 16640
rect 30561 16609 30573 16612
rect 30607 16609 30619 16643
rect 34698 16640 34704 16652
rect 30561 16603 30619 16609
rect 34440 16612 34704 16640
rect 30101 16575 30159 16581
rect 30101 16541 30113 16575
rect 30147 16541 30159 16575
rect 30101 16535 30159 16541
rect 30469 16575 30527 16581
rect 30469 16541 30481 16575
rect 30515 16541 30527 16575
rect 30469 16535 30527 16541
rect 27764 16476 28948 16504
rect 27764 16464 27770 16476
rect 29638 16464 29644 16516
rect 29696 16504 29702 16516
rect 30374 16504 30380 16516
rect 29696 16476 30380 16504
rect 29696 16464 29702 16476
rect 30374 16464 30380 16476
rect 30432 16504 30438 16516
rect 30484 16504 30512 16535
rect 30926 16532 30932 16584
rect 30984 16572 30990 16584
rect 31205 16575 31263 16581
rect 31205 16572 31217 16575
rect 30984 16544 31217 16572
rect 30984 16532 30990 16544
rect 31205 16541 31217 16544
rect 31251 16541 31263 16575
rect 31478 16572 31484 16584
rect 31439 16544 31484 16572
rect 31205 16535 31263 16541
rect 31478 16532 31484 16544
rect 31536 16532 31542 16584
rect 32766 16572 32772 16584
rect 31726 16544 32444 16572
rect 32727 16544 32772 16572
rect 30432 16476 30512 16504
rect 30432 16464 30438 16476
rect 31018 16464 31024 16516
rect 31076 16504 31082 16516
rect 31297 16507 31355 16513
rect 31297 16504 31309 16507
rect 31076 16476 31309 16504
rect 31076 16464 31082 16476
rect 31297 16473 31309 16476
rect 31343 16504 31355 16507
rect 31726 16504 31754 16544
rect 31343 16476 31754 16504
rect 31343 16473 31355 16476
rect 31297 16467 31355 16473
rect 32214 16464 32220 16516
rect 32272 16504 32278 16516
rect 32309 16507 32367 16513
rect 32309 16504 32321 16507
rect 32272 16476 32321 16504
rect 32272 16464 32278 16476
rect 32309 16473 32321 16476
rect 32355 16473 32367 16507
rect 32416 16504 32444 16544
rect 32766 16532 32772 16544
rect 32824 16532 32830 16584
rect 33042 16572 33048 16584
rect 33003 16544 33048 16572
rect 33042 16532 33048 16544
rect 33100 16572 33106 16584
rect 34440 16572 34468 16612
rect 34698 16600 34704 16612
rect 34756 16640 34762 16652
rect 34977 16643 35035 16649
rect 34977 16640 34989 16643
rect 34756 16612 34989 16640
rect 34756 16600 34762 16612
rect 34977 16609 34989 16612
rect 35023 16609 35035 16643
rect 34977 16603 35035 16609
rect 35342 16600 35348 16652
rect 35400 16640 35406 16652
rect 35400 16612 35664 16640
rect 35400 16600 35406 16612
rect 33100 16544 34468 16572
rect 33100 16532 33106 16544
rect 34514 16532 34520 16584
rect 34572 16572 34578 16584
rect 35636 16581 35664 16612
rect 35894 16600 35900 16652
rect 35952 16640 35958 16652
rect 36265 16643 36323 16649
rect 36265 16640 36277 16643
rect 35952 16612 36277 16640
rect 35952 16600 35958 16612
rect 36265 16609 36277 16612
rect 36311 16609 36323 16643
rect 36265 16603 36323 16609
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 34572 16544 34897 16572
rect 34572 16532 34578 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 35621 16575 35679 16581
rect 35621 16541 35633 16575
rect 35667 16541 35679 16575
rect 35621 16535 35679 16541
rect 32861 16507 32919 16513
rect 32861 16504 32873 16507
rect 32416 16476 32873 16504
rect 32309 16467 32367 16473
rect 32861 16473 32873 16476
rect 32907 16504 32919 16507
rect 33318 16504 33324 16516
rect 32907 16476 33324 16504
rect 32907 16473 32919 16476
rect 32861 16467 32919 16473
rect 33318 16464 33324 16476
rect 33376 16464 33382 16516
rect 33686 16504 33692 16516
rect 33647 16476 33692 16504
rect 33686 16464 33692 16476
rect 33744 16464 33750 16516
rect 35161 16507 35219 16513
rect 35161 16473 35173 16507
rect 35207 16504 35219 16507
rect 36262 16504 36268 16516
rect 35207 16476 36268 16504
rect 35207 16473 35219 16476
rect 35161 16467 35219 16473
rect 36262 16464 36268 16476
rect 36320 16464 36326 16516
rect 36449 16507 36507 16513
rect 36449 16473 36461 16507
rect 36495 16504 36507 16507
rect 37918 16504 37924 16516
rect 36495 16476 37924 16504
rect 36495 16473 36507 16476
rect 36449 16467 36507 16473
rect 37918 16464 37924 16476
rect 37976 16464 37982 16516
rect 38102 16504 38108 16516
rect 38063 16476 38108 16504
rect 38102 16464 38108 16476
rect 38160 16464 38166 16516
rect 23348 16408 23520 16436
rect 23348 16396 23354 16408
rect 24854 16396 24860 16448
rect 24912 16396 24918 16448
rect 25317 16439 25375 16445
rect 25317 16405 25329 16439
rect 25363 16436 25375 16439
rect 25498 16436 25504 16448
rect 25363 16408 25504 16436
rect 25363 16405 25375 16408
rect 25317 16399 25375 16405
rect 25498 16396 25504 16408
rect 25556 16436 25562 16448
rect 25774 16436 25780 16448
rect 25556 16408 25780 16436
rect 25556 16396 25562 16408
rect 25774 16396 25780 16408
rect 25832 16396 25838 16448
rect 25961 16439 26019 16445
rect 25961 16405 25973 16439
rect 26007 16436 26019 16439
rect 28074 16436 28080 16448
rect 26007 16408 28080 16436
rect 26007 16405 26019 16408
rect 25961 16399 26019 16405
rect 28074 16396 28080 16408
rect 28132 16396 28138 16448
rect 28169 16439 28227 16445
rect 28169 16405 28181 16439
rect 28215 16436 28227 16439
rect 28258 16436 28264 16448
rect 28215 16408 28264 16436
rect 28215 16405 28227 16408
rect 28169 16399 28227 16405
rect 28258 16396 28264 16408
rect 28316 16396 28322 16448
rect 29730 16396 29736 16448
rect 29788 16436 29794 16448
rect 30098 16436 30104 16448
rect 29788 16408 30104 16436
rect 29788 16396 29794 16408
rect 30098 16396 30104 16408
rect 30156 16436 30162 16448
rect 30193 16439 30251 16445
rect 30193 16436 30205 16439
rect 30156 16408 30205 16436
rect 30156 16396 30162 16408
rect 30193 16405 30205 16408
rect 30239 16405 30251 16439
rect 30193 16399 30251 16405
rect 30285 16439 30343 16445
rect 30285 16405 30297 16439
rect 30331 16436 30343 16439
rect 30466 16436 30472 16448
rect 30331 16408 30472 16436
rect 30331 16405 30343 16408
rect 30285 16399 30343 16405
rect 30466 16396 30472 16408
rect 30524 16396 30530 16448
rect 30742 16436 30748 16448
rect 30703 16408 30748 16436
rect 30742 16396 30748 16408
rect 30800 16396 30806 16448
rect 32109 16439 32167 16445
rect 32109 16405 32121 16439
rect 32155 16436 32167 16439
rect 32490 16436 32496 16448
rect 32155 16408 32496 16436
rect 32155 16405 32167 16408
rect 32109 16399 32167 16405
rect 32490 16396 32496 16408
rect 32548 16396 32554 16448
rect 33229 16439 33287 16445
rect 33229 16405 33241 16439
rect 33275 16436 33287 16439
rect 33889 16439 33947 16445
rect 33889 16436 33901 16439
rect 33275 16408 33901 16436
rect 33275 16405 33287 16408
rect 33229 16399 33287 16405
rect 33889 16405 33901 16408
rect 33935 16405 33947 16439
rect 33889 16399 33947 16405
rect 34790 16396 34796 16448
rect 34848 16436 34854 16448
rect 35713 16439 35771 16445
rect 35713 16436 35725 16439
rect 34848 16408 35725 16436
rect 34848 16396 34854 16408
rect 35713 16405 35725 16408
rect 35759 16405 35771 16439
rect 35713 16399 35771 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 9214 16232 9220 16244
rect 9175 16204 9220 16232
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 12894 16232 12900 16244
rect 12855 16204 12900 16232
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 14182 16192 14188 16244
rect 14240 16232 14246 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14240 16204 15025 16232
rect 14240 16192 14246 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 15013 16195 15071 16201
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20438 16192 20444 16244
rect 20496 16232 20502 16244
rect 23014 16232 23020 16244
rect 20496 16204 23020 16232
rect 20496 16192 20502 16204
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 23293 16235 23351 16241
rect 23293 16201 23305 16235
rect 23339 16232 23351 16235
rect 27614 16232 27620 16244
rect 23339 16204 27620 16232
rect 23339 16201 23351 16204
rect 23293 16195 23351 16201
rect 27614 16192 27620 16204
rect 27672 16192 27678 16244
rect 29638 16232 29644 16244
rect 29599 16204 29644 16232
rect 29638 16192 29644 16204
rect 29696 16192 29702 16244
rect 30101 16235 30159 16241
rect 30101 16201 30113 16235
rect 30147 16232 30159 16235
rect 31110 16232 31116 16244
rect 30147 16204 31116 16232
rect 30147 16201 30159 16204
rect 30101 16195 30159 16201
rect 31110 16192 31116 16204
rect 31168 16192 31174 16244
rect 32769 16235 32827 16241
rect 32769 16201 32781 16235
rect 32815 16232 32827 16235
rect 34790 16232 34796 16244
rect 32815 16204 34796 16232
rect 32815 16201 32827 16204
rect 32769 16195 32827 16201
rect 34790 16192 34796 16204
rect 34848 16192 34854 16244
rect 37277 16235 37335 16241
rect 37277 16232 37289 16235
rect 36280 16204 37289 16232
rect 8662 16124 8668 16176
rect 8720 16164 8726 16176
rect 10689 16167 10747 16173
rect 10689 16164 10701 16167
rect 8720 16136 10701 16164
rect 8720 16124 8726 16136
rect 10689 16133 10701 16136
rect 10735 16133 10747 16167
rect 10689 16127 10747 16133
rect 10873 16167 10931 16173
rect 10873 16133 10885 16167
rect 10919 16164 10931 16167
rect 12618 16164 12624 16176
rect 10919 16136 12624 16164
rect 10919 16133 10931 16136
rect 10873 16127 10931 16133
rect 12618 16124 12624 16136
rect 12676 16124 12682 16176
rect 14734 16164 14740 16176
rect 13648 16136 14740 16164
rect 9398 16096 9404 16108
rect 9359 16068 9404 16096
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 13648 16105 13676 16136
rect 14734 16124 14740 16136
rect 14792 16124 14798 16176
rect 18138 16124 18144 16176
rect 18196 16164 18202 16176
rect 18196 16136 18722 16164
rect 18196 16124 18202 16136
rect 20622 16124 20628 16176
rect 20680 16164 20686 16176
rect 20680 16136 22094 16164
rect 20680 16124 20686 16136
rect 13906 16105 13912 16108
rect 11773 16099 11831 16105
rect 11773 16096 11785 16099
rect 11020 16068 11785 16096
rect 11020 16056 11026 16068
rect 11773 16065 11785 16068
rect 11819 16065 11831 16099
rect 11773 16059 11831 16065
rect 13633 16099 13691 16105
rect 13633 16065 13645 16099
rect 13679 16065 13691 16099
rect 13900 16096 13912 16105
rect 13867 16068 13912 16096
rect 13633 16059 13691 16065
rect 13900 16059 13912 16068
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 2133 15895 2191 15901
rect 2133 15861 2145 15895
rect 2179 15892 2191 15895
rect 3234 15892 3240 15904
rect 2179 15864 3240 15892
rect 2179 15861 2191 15864
rect 2133 15855 2191 15861
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 11532 15892 11560 15991
rect 13648 15960 13676 16059
rect 13906 16056 13912 16059
rect 13964 16056 13970 16108
rect 15746 16096 15752 16108
rect 15707 16068 15752 16096
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 17126 16096 17132 16108
rect 17087 16068 17132 16096
rect 17126 16056 17132 16068
rect 17184 16056 17190 16108
rect 20346 16096 20352 16108
rect 20307 16068 20352 16096
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 21082 16096 21088 16108
rect 21043 16068 21088 16096
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 22066 16096 22094 16136
rect 23198 16124 23204 16176
rect 23256 16164 23262 16176
rect 23845 16167 23903 16173
rect 23845 16164 23857 16167
rect 23256 16136 23857 16164
rect 23256 16124 23262 16136
rect 23845 16133 23857 16136
rect 23891 16164 23903 16167
rect 24854 16164 24860 16176
rect 23891 16136 24860 16164
rect 23891 16133 23903 16136
rect 23845 16127 23903 16133
rect 24854 16124 24860 16136
rect 24912 16124 24918 16176
rect 25038 16124 25044 16176
rect 25096 16164 25102 16176
rect 25096 16136 27752 16164
rect 25096 16124 25102 16136
rect 22186 16096 22192 16108
rect 22066 16068 22192 16096
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22370 16096 22376 16108
rect 22331 16068 22376 16096
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 23106 16096 23112 16108
rect 23067 16068 23112 16096
rect 23106 16056 23112 16068
rect 23164 16056 23170 16108
rect 24210 16096 24216 16108
rect 24171 16068 24216 16096
rect 24210 16056 24216 16068
rect 24268 16056 24274 16108
rect 24946 16096 24952 16108
rect 24907 16068 24952 16096
rect 24946 16056 24952 16068
rect 25004 16056 25010 16108
rect 25774 16096 25780 16108
rect 25735 16068 25780 16096
rect 25774 16056 25780 16068
rect 25832 16056 25838 16108
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16096 26111 16099
rect 26694 16096 26700 16108
rect 26099 16068 26700 16096
rect 26099 16065 26111 16068
rect 26053 16059 26111 16065
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 27154 16096 27160 16108
rect 27115 16068 27160 16096
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27246 16056 27252 16108
rect 27304 16096 27310 16108
rect 27341 16099 27399 16105
rect 27341 16096 27353 16099
rect 27304 16068 27353 16096
rect 27304 16056 27310 16068
rect 27341 16065 27353 16068
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 27433 16099 27491 16105
rect 27433 16065 27445 16099
rect 27479 16096 27491 16099
rect 27614 16096 27620 16108
rect 27479 16068 27620 16096
rect 27479 16065 27491 16068
rect 27433 16059 27491 16065
rect 27614 16056 27620 16068
rect 27672 16056 27678 16108
rect 27724 16096 27752 16136
rect 28074 16124 28080 16176
rect 28132 16164 28138 16176
rect 32677 16167 32735 16173
rect 28132 16136 28658 16164
rect 28132 16124 28138 16136
rect 32677 16133 32689 16167
rect 32723 16164 32735 16167
rect 33134 16164 33140 16176
rect 32723 16136 33140 16164
rect 32723 16133 32735 16136
rect 32677 16127 32735 16133
rect 33134 16124 33140 16136
rect 33192 16164 33198 16176
rect 33870 16164 33876 16176
rect 33192 16136 33876 16164
rect 33192 16124 33198 16136
rect 33870 16124 33876 16136
rect 33928 16124 33934 16176
rect 34149 16167 34207 16173
rect 34149 16133 34161 16167
rect 34195 16164 34207 16167
rect 34514 16164 34520 16176
rect 34195 16136 34520 16164
rect 34195 16133 34207 16136
rect 34149 16127 34207 16133
rect 34514 16124 34520 16136
rect 34572 16124 34578 16176
rect 35526 16124 35532 16176
rect 35584 16124 35590 16176
rect 36280 16173 36308 16204
rect 37277 16201 37289 16204
rect 37323 16201 37335 16235
rect 37277 16195 37335 16201
rect 37918 16192 37924 16244
rect 37976 16232 37982 16244
rect 38013 16235 38071 16241
rect 38013 16232 38025 16235
rect 37976 16204 38025 16232
rect 37976 16192 37982 16204
rect 38013 16201 38025 16204
rect 38059 16201 38071 16235
rect 38013 16195 38071 16201
rect 36265 16167 36323 16173
rect 36265 16133 36277 16167
rect 36311 16133 36323 16167
rect 36265 16127 36323 16133
rect 27893 16099 27951 16105
rect 27893 16096 27905 16099
rect 27724 16068 27905 16096
rect 27893 16065 27905 16068
rect 27939 16065 27951 16099
rect 27893 16059 27951 16065
rect 30469 16099 30527 16105
rect 30469 16065 30481 16099
rect 30515 16096 30527 16099
rect 30742 16096 30748 16108
rect 30515 16068 30748 16096
rect 30515 16065 30527 16068
rect 30469 16059 30527 16065
rect 30742 16056 30748 16068
rect 30800 16056 30806 16108
rect 31386 16096 31392 16108
rect 31347 16068 31392 16096
rect 31386 16056 31392 16068
rect 31444 16056 31450 16108
rect 32950 16056 32956 16108
rect 33008 16096 33014 16108
rect 34054 16096 34060 16108
rect 33008 16068 34060 16096
rect 33008 16056 33014 16068
rect 34054 16056 34060 16068
rect 34112 16056 34118 16108
rect 34333 16099 34391 16105
rect 34333 16065 34345 16099
rect 34379 16096 34391 16099
rect 34790 16096 34796 16108
rect 34379 16068 34796 16096
rect 34379 16065 34391 16068
rect 34333 16059 34391 16065
rect 34790 16056 34796 16068
rect 34848 16056 34854 16108
rect 37458 16096 37464 16108
rect 37419 16068 37464 16096
rect 37458 16056 37464 16068
rect 37516 16056 37522 16108
rect 37826 16056 37832 16108
rect 37884 16096 37890 16108
rect 37921 16099 37979 16105
rect 37921 16096 37933 16099
rect 37884 16068 37933 16096
rect 37884 16056 37890 16068
rect 37921 16065 37933 16068
rect 37967 16065 37979 16099
rect 37921 16059 37979 16065
rect 17862 16028 17868 16040
rect 12820 15932 13676 15960
rect 17236 16000 17868 16028
rect 12710 15892 12716 15904
rect 11532 15864 12716 15892
rect 12710 15852 12716 15864
rect 12768 15892 12774 15904
rect 12820 15892 12848 15932
rect 15838 15892 15844 15904
rect 12768 15864 12848 15892
rect 15799 15864 15844 15892
rect 12768 15852 12774 15864
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 17236 15901 17264 16000
rect 17862 15988 17868 16000
rect 17920 16028 17926 16040
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 17920 16000 17969 16028
rect 17920 15988 17926 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 18230 16028 18236 16040
rect 18191 16000 18236 16028
rect 17957 15991 18015 15997
rect 18230 15988 18236 16000
rect 18288 15988 18294 16040
rect 22833 16031 22891 16037
rect 22833 15997 22845 16031
rect 22879 16028 22891 16031
rect 24486 16028 24492 16040
rect 22879 16000 24492 16028
rect 22879 15997 22891 16000
rect 22833 15991 22891 15997
rect 20530 15920 20536 15972
rect 20588 15960 20594 15972
rect 22848 15960 22876 15991
rect 24486 15988 24492 16000
rect 24544 15988 24550 16040
rect 25961 16031 26019 16037
rect 25961 15997 25973 16031
rect 26007 16028 26019 16031
rect 30282 16028 30288 16040
rect 26007 16000 30288 16028
rect 26007 15997 26019 16000
rect 25961 15991 26019 15997
rect 30282 15988 30288 16000
rect 30340 15988 30346 16040
rect 30377 16031 30435 16037
rect 30377 15997 30389 16031
rect 30423 16028 30435 16031
rect 30423 16000 31754 16028
rect 30423 15997 30435 16000
rect 30377 15991 30435 15997
rect 20588 15932 22876 15960
rect 25041 15963 25099 15969
rect 20588 15920 20594 15932
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 16724 15864 17233 15892
rect 16724 15852 16730 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 19705 15895 19763 15901
rect 19705 15861 19717 15895
rect 19751 15892 19763 15895
rect 19794 15892 19800 15904
rect 19751 15864 19800 15892
rect 19751 15861 19763 15864
rect 19705 15855 19763 15861
rect 19794 15852 19800 15864
rect 19852 15852 19858 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21542 15892 21548 15904
rect 21315 15864 21548 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 22112 15901 22140 15932
rect 25041 15929 25053 15963
rect 25087 15960 25099 15963
rect 27430 15960 27436 15972
rect 25087 15932 27436 15960
rect 25087 15929 25099 15932
rect 25041 15923 25099 15929
rect 27430 15920 27436 15932
rect 27488 15920 27494 15972
rect 29178 15920 29184 15972
rect 29236 15960 29242 15972
rect 30466 15960 30472 15972
rect 29236 15932 30472 15960
rect 29236 15920 29242 15932
rect 30466 15920 30472 15932
rect 30524 15920 30530 15972
rect 31726 15960 31754 16000
rect 32582 15988 32588 16040
rect 32640 16028 32646 16040
rect 33045 16031 33103 16037
rect 33045 16028 33057 16031
rect 32640 16000 33057 16028
rect 32640 15988 32646 16000
rect 33045 15997 33057 16000
rect 33091 15997 33103 16031
rect 36538 16028 36544 16040
rect 36499 16000 36544 16028
rect 33045 15991 33103 15997
rect 36538 15988 36544 16000
rect 36596 15988 36602 16040
rect 31726 15932 34468 15960
rect 22097 15895 22155 15901
rect 22097 15861 22109 15895
rect 22143 15892 22155 15895
rect 22922 15892 22928 15904
rect 22143 15864 22177 15892
rect 22883 15864 22928 15892
rect 22143 15861 22155 15864
rect 22097 15855 22155 15861
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 25498 15852 25504 15904
rect 25556 15892 25562 15904
rect 25593 15895 25651 15901
rect 25593 15892 25605 15895
rect 25556 15864 25605 15892
rect 25556 15852 25562 15864
rect 25593 15861 25605 15864
rect 25639 15861 25651 15895
rect 25593 15855 25651 15861
rect 27157 15895 27215 15901
rect 27157 15861 27169 15895
rect 27203 15892 27215 15895
rect 27982 15892 27988 15904
rect 27203 15864 27988 15892
rect 27203 15861 27215 15864
rect 27157 15855 27215 15861
rect 27982 15852 27988 15864
rect 28040 15852 28046 15904
rect 28156 15895 28214 15901
rect 28156 15861 28168 15895
rect 28202 15892 28214 15895
rect 28350 15892 28356 15904
rect 28202 15864 28356 15892
rect 28202 15861 28214 15864
rect 28156 15855 28214 15861
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 31481 15895 31539 15901
rect 31481 15861 31493 15895
rect 31527 15892 31539 15895
rect 31662 15892 31668 15904
rect 31527 15864 31668 15892
rect 31527 15861 31539 15864
rect 31481 15855 31539 15861
rect 31662 15852 31668 15864
rect 31720 15852 31726 15904
rect 32950 15892 32956 15904
rect 32911 15864 32956 15892
rect 32950 15852 32956 15864
rect 33008 15852 33014 15904
rect 33137 15895 33195 15901
rect 33137 15861 33149 15895
rect 33183 15892 33195 15895
rect 33318 15892 33324 15904
rect 33183 15864 33324 15892
rect 33183 15861 33195 15864
rect 33137 15855 33195 15861
rect 33318 15852 33324 15864
rect 33376 15852 33382 15904
rect 34330 15892 34336 15904
rect 34291 15864 34336 15892
rect 34330 15852 34336 15864
rect 34388 15852 34394 15904
rect 34440 15892 34468 15932
rect 34698 15920 34704 15972
rect 34756 15960 34762 15972
rect 34793 15963 34851 15969
rect 34793 15960 34805 15963
rect 34756 15932 34805 15960
rect 34756 15920 34762 15932
rect 34793 15929 34805 15932
rect 34839 15929 34851 15963
rect 34793 15923 34851 15929
rect 35710 15892 35716 15904
rect 34440 15864 35716 15892
rect 35710 15852 35716 15864
rect 35768 15852 35774 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 10962 15688 10968 15700
rect 10923 15660 10968 15688
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 13136 15660 13553 15688
rect 13136 15648 13142 15660
rect 13541 15657 13553 15660
rect 13587 15688 13599 15691
rect 13630 15688 13636 15700
rect 13587 15660 13636 15688
rect 13587 15657 13599 15660
rect 13541 15651 13599 15657
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 18230 15648 18236 15700
rect 18288 15688 18294 15700
rect 18417 15691 18475 15697
rect 18417 15688 18429 15691
rect 18288 15660 18429 15688
rect 18288 15648 18294 15660
rect 18417 15657 18429 15660
rect 18463 15657 18475 15691
rect 18417 15651 18475 15657
rect 18874 15648 18880 15700
rect 18932 15688 18938 15700
rect 20625 15691 20683 15697
rect 20625 15688 20637 15691
rect 18932 15660 20637 15688
rect 18932 15648 18938 15660
rect 20625 15657 20637 15660
rect 20671 15657 20683 15691
rect 20625 15651 20683 15657
rect 24673 15691 24731 15697
rect 24673 15657 24685 15691
rect 24719 15688 24731 15691
rect 28074 15688 28080 15700
rect 24719 15660 28080 15688
rect 24719 15657 24731 15660
rect 24673 15651 24731 15657
rect 28074 15648 28080 15660
rect 28132 15648 28138 15700
rect 28350 15648 28356 15700
rect 28408 15688 28414 15700
rect 28445 15691 28503 15697
rect 28445 15688 28457 15691
rect 28408 15660 28457 15688
rect 28408 15648 28414 15660
rect 28445 15657 28457 15660
rect 28491 15657 28503 15691
rect 28445 15651 28503 15657
rect 29641 15691 29699 15697
rect 29641 15657 29653 15691
rect 29687 15688 29699 15691
rect 33134 15688 33140 15700
rect 29687 15660 33140 15688
rect 29687 15657 29699 15660
rect 29641 15651 29699 15657
rect 33134 15648 33140 15660
rect 33192 15648 33198 15700
rect 34790 15648 34796 15700
rect 34848 15688 34854 15700
rect 35345 15691 35403 15697
rect 35345 15688 35357 15691
rect 34848 15660 35357 15688
rect 34848 15648 34854 15660
rect 35345 15657 35357 15660
rect 35391 15657 35403 15691
rect 35345 15651 35403 15657
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 10008 15592 11529 15620
rect 10008 15580 10014 15592
rect 11517 15589 11529 15592
rect 11563 15589 11575 15623
rect 11517 15583 11575 15589
rect 13906 15580 13912 15632
rect 13964 15620 13970 15632
rect 14369 15623 14427 15629
rect 14369 15620 14381 15623
rect 13964 15592 14381 15620
rect 13964 15580 13970 15592
rect 14369 15589 14381 15592
rect 14415 15620 14427 15623
rect 14734 15620 14740 15632
rect 14415 15592 14740 15620
rect 14415 15589 14427 15592
rect 14369 15583 14427 15589
rect 14734 15580 14740 15592
rect 14792 15580 14798 15632
rect 19245 15623 19303 15629
rect 19245 15589 19257 15623
rect 19291 15589 19303 15623
rect 19245 15583 19303 15589
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 3234 15552 3240 15564
rect 3195 15524 3240 15552
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 14752 15552 14780 15580
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 14752 15524 14841 15552
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 16623 15524 17908 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 17880 15496 17908 15524
rect 10778 15484 10784 15496
rect 10739 15456 10784 15484
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 11422 15484 11428 15496
rect 11383 15456 11428 15484
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15484 11667 15487
rect 11882 15484 11888 15496
rect 11655 15456 11888 15484
rect 11655 15453 11667 15456
rect 11609 15447 11667 15453
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15484 12219 15487
rect 12710 15484 12716 15496
rect 12207 15456 12716 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 17678 15484 17684 15496
rect 17639 15456 17684 15484
rect 17678 15444 17684 15456
rect 17736 15444 17742 15496
rect 17862 15484 17868 15496
rect 17823 15456 17868 15484
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 19260 15484 19288 15583
rect 20438 15580 20444 15632
rect 20496 15620 20502 15632
rect 22002 15620 22008 15632
rect 20496 15592 22008 15620
rect 20496 15580 20502 15592
rect 22002 15580 22008 15592
rect 22060 15580 22066 15632
rect 22554 15580 22560 15632
rect 22612 15620 22618 15632
rect 22741 15623 22799 15629
rect 22741 15620 22753 15623
rect 22612 15592 22753 15620
rect 22612 15580 22618 15592
rect 22741 15589 22753 15592
rect 22787 15620 22799 15623
rect 23198 15620 23204 15632
rect 22787 15592 23204 15620
rect 22787 15589 22799 15592
rect 22741 15583 22799 15589
rect 23198 15580 23204 15592
rect 23256 15580 23262 15632
rect 26694 15580 26700 15632
rect 26752 15620 26758 15632
rect 26973 15623 27031 15629
rect 26973 15620 26985 15623
rect 26752 15592 26985 15620
rect 26752 15580 26758 15592
rect 26973 15589 26985 15592
rect 27019 15589 27031 15623
rect 32306 15620 32312 15632
rect 26973 15583 27031 15589
rect 29564 15592 32312 15620
rect 19794 15552 19800 15564
rect 19755 15524 19800 15552
rect 19794 15512 19800 15524
rect 19852 15552 19858 15564
rect 20809 15555 20867 15561
rect 19852 15524 20668 15552
rect 19852 15512 19858 15524
rect 20640 15493 20668 15524
rect 20809 15521 20821 15555
rect 20855 15552 20867 15555
rect 21082 15552 21088 15564
rect 20855 15524 21088 15552
rect 20855 15521 20867 15524
rect 20809 15515 20867 15521
rect 21082 15512 21088 15524
rect 21140 15512 21146 15564
rect 25038 15512 25044 15564
rect 25096 15552 25102 15564
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 25096 15524 25237 15552
rect 25096 15512 25102 15524
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25498 15552 25504 15564
rect 25459 15524 25504 15552
rect 25225 15515 25283 15521
rect 25498 15512 25504 15524
rect 25556 15512 25562 15564
rect 27982 15552 27988 15564
rect 27943 15524 27988 15552
rect 27982 15512 27988 15524
rect 28040 15512 28046 15564
rect 18647 15456 19288 15484
rect 20625 15487 20683 15493
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20898 15484 20904 15496
rect 20859 15456 20904 15484
rect 20625 15447 20683 15453
rect 20898 15444 20904 15456
rect 20956 15484 20962 15496
rect 21818 15484 21824 15496
rect 20956 15456 21824 15484
rect 20956 15444 20962 15456
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22244 15456 22569 15484
rect 22244 15444 22250 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15484 23903 15487
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 23891 15456 24593 15484
rect 23891 15453 23903 15456
rect 23845 15447 23903 15453
rect 24581 15453 24593 15456
rect 24627 15484 24639 15487
rect 24946 15484 24952 15496
rect 24627 15456 24952 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 27798 15444 27804 15496
rect 27856 15484 27862 15496
rect 28077 15487 28135 15493
rect 28077 15484 28089 15487
rect 27856 15456 28089 15484
rect 27856 15444 27862 15456
rect 28077 15453 28089 15456
rect 28123 15453 28135 15487
rect 28258 15484 28264 15496
rect 28219 15456 28264 15484
rect 28077 15447 28135 15453
rect 28258 15444 28264 15456
rect 28316 15444 28322 15496
rect 29564 15493 29592 15592
rect 32306 15580 32312 15592
rect 32364 15580 32370 15632
rect 30190 15552 30196 15564
rect 30151 15524 30196 15552
rect 30190 15512 30196 15524
rect 30248 15512 30254 15564
rect 31573 15555 31631 15561
rect 31573 15552 31585 15555
rect 31220 15524 31585 15552
rect 31220 15496 31248 15524
rect 31573 15521 31585 15524
rect 31619 15521 31631 15555
rect 31573 15515 31631 15521
rect 31662 15512 31668 15564
rect 31720 15552 31726 15564
rect 32401 15555 32459 15561
rect 32401 15552 32413 15555
rect 31720 15524 32413 15552
rect 31720 15512 31726 15524
rect 32401 15521 32413 15524
rect 32447 15521 32459 15555
rect 32401 15515 32459 15521
rect 32677 15555 32735 15561
rect 32677 15521 32689 15555
rect 32723 15552 32735 15555
rect 34330 15552 34336 15564
rect 32723 15524 34336 15552
rect 32723 15521 32735 15524
rect 32677 15515 32735 15521
rect 34330 15512 34336 15524
rect 34388 15512 34394 15564
rect 35250 15552 35256 15564
rect 35211 15524 35256 15552
rect 35250 15512 35256 15524
rect 35308 15512 35314 15564
rect 37090 15552 37096 15564
rect 37051 15524 37096 15552
rect 37090 15512 37096 15524
rect 37148 15512 37154 15564
rect 29549 15487 29607 15493
rect 29549 15453 29561 15487
rect 29595 15453 29607 15487
rect 29730 15484 29736 15496
rect 29691 15456 29736 15484
rect 29549 15447 29607 15453
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 30374 15484 30380 15496
rect 30335 15456 30380 15484
rect 30374 15444 30380 15456
rect 30432 15444 30438 15496
rect 30466 15444 30472 15496
rect 30524 15484 30530 15496
rect 30745 15487 30803 15493
rect 30524 15456 30569 15484
rect 30524 15444 30530 15456
rect 30745 15453 30757 15487
rect 30791 15484 30803 15487
rect 31202 15484 31208 15496
rect 30791 15456 31208 15484
rect 30791 15453 30803 15456
rect 30745 15447 30803 15453
rect 31202 15444 31208 15456
rect 31260 15444 31266 15496
rect 31389 15487 31447 15493
rect 31389 15453 31401 15487
rect 31435 15484 31447 15487
rect 31478 15484 31484 15496
rect 31435 15456 31484 15484
rect 31435 15453 31447 15456
rect 31389 15447 31447 15453
rect 31478 15444 31484 15456
rect 31536 15444 31542 15496
rect 34054 15444 34060 15496
rect 34112 15484 34118 15496
rect 35434 15484 35440 15496
rect 34112 15456 35440 15484
rect 34112 15444 34118 15456
rect 35434 15444 35440 15456
rect 35492 15444 35498 15496
rect 35529 15487 35587 15493
rect 35529 15453 35541 15487
rect 35575 15484 35587 15487
rect 35618 15484 35624 15496
rect 35575 15456 35624 15484
rect 35575 15453 35587 15456
rect 35529 15447 35587 15453
rect 35618 15444 35624 15456
rect 35676 15444 35682 15496
rect 38102 15444 38108 15496
rect 38160 15484 38166 15496
rect 38160 15456 38205 15484
rect 38160 15444 38166 15456
rect 3050 15416 3056 15428
rect 3011 15388 3056 15416
rect 3050 15376 3056 15388
rect 3108 15376 3114 15428
rect 12428 15419 12486 15425
rect 12428 15385 12440 15419
rect 12474 15416 12486 15419
rect 12526 15416 12532 15428
rect 12474 15388 12532 15416
rect 12474 15385 12486 15388
rect 12428 15379 12486 15385
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 12618 15376 12624 15428
rect 12676 15416 12682 15428
rect 14185 15419 14243 15425
rect 14185 15416 14197 15419
rect 12676 15388 14197 15416
rect 12676 15376 12682 15388
rect 14185 15385 14197 15388
rect 14231 15385 14243 15419
rect 15102 15416 15108 15428
rect 15063 15388 15108 15416
rect 14185 15379 14243 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 15838 15376 15844 15428
rect 15896 15376 15902 15428
rect 21542 15416 21548 15428
rect 21503 15388 21548 15416
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 21729 15419 21787 15425
rect 21729 15385 21741 15419
rect 21775 15416 21787 15419
rect 22002 15416 22008 15428
rect 21775 15388 22008 15416
rect 21775 15385 21787 15388
rect 21729 15379 21787 15385
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 23753 15419 23811 15425
rect 23753 15385 23765 15419
rect 23799 15416 23811 15419
rect 34698 15416 34704 15428
rect 23799 15388 25990 15416
rect 30484 15388 31248 15416
rect 33902 15388 34704 15416
rect 23799 15385 23811 15388
rect 23753 15379 23811 15385
rect 17494 15348 17500 15360
rect 17455 15320 17500 15348
rect 17494 15308 17500 15320
rect 17552 15308 17558 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 19484 15320 19625 15348
rect 19484 15308 19490 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 19705 15351 19763 15357
rect 19705 15317 19717 15351
rect 19751 15348 19763 15351
rect 19978 15348 19984 15360
rect 19751 15320 19984 15348
rect 19751 15317 19763 15320
rect 19705 15311 19763 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20441 15351 20499 15357
rect 20441 15317 20453 15351
rect 20487 15348 20499 15351
rect 20530 15348 20536 15360
rect 20487 15320 20536 15348
rect 20487 15317 20499 15320
rect 20441 15311 20499 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 20898 15308 20904 15360
rect 20956 15348 20962 15360
rect 21361 15351 21419 15357
rect 21361 15348 21373 15351
rect 20956 15320 21373 15348
rect 20956 15308 20962 15320
rect 21361 15317 21373 15320
rect 21407 15317 21419 15351
rect 21361 15311 21419 15317
rect 26418 15308 26424 15360
rect 26476 15348 26482 15360
rect 26878 15348 26884 15360
rect 26476 15320 26884 15348
rect 26476 15308 26482 15320
rect 26878 15308 26884 15320
rect 26936 15348 26942 15360
rect 30484 15348 30512 15388
rect 26936 15320 30512 15348
rect 26936 15308 26942 15320
rect 30558 15308 30564 15360
rect 30616 15348 30622 15360
rect 31220 15357 31248 15388
rect 34698 15376 34704 15388
rect 34756 15376 34762 15428
rect 37918 15416 37924 15428
rect 37879 15388 37924 15416
rect 37918 15376 37924 15388
rect 37976 15376 37982 15428
rect 31205 15351 31263 15357
rect 30616 15320 30661 15348
rect 30616 15308 30622 15320
rect 31205 15317 31217 15351
rect 31251 15317 31263 15351
rect 31205 15311 31263 15317
rect 34149 15351 34207 15357
rect 34149 15317 34161 15351
rect 34195 15348 34207 15351
rect 34514 15348 34520 15360
rect 34195 15320 34520 15348
rect 34195 15317 34207 15320
rect 34149 15311 34207 15317
rect 34514 15308 34520 15320
rect 34572 15348 34578 15360
rect 34790 15348 34796 15360
rect 34572 15320 34796 15348
rect 34572 15308 34578 15320
rect 34790 15308 34796 15320
rect 34848 15308 34854 15360
rect 35250 15308 35256 15360
rect 35308 15348 35314 15360
rect 35710 15348 35716 15360
rect 35308 15320 35716 15348
rect 35308 15308 35314 15320
rect 35710 15308 35716 15320
rect 35768 15308 35774 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 2685 15147 2743 15153
rect 2685 15113 2697 15147
rect 2731 15144 2743 15147
rect 3050 15144 3056 15156
rect 2731 15116 3056 15144
rect 2731 15113 2743 15116
rect 2685 15107 2743 15113
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 13817 15147 13875 15153
rect 13817 15113 13829 15147
rect 13863 15144 13875 15147
rect 14458 15144 14464 15156
rect 13863 15116 14464 15144
rect 13863 15113 13875 15116
rect 13817 15107 13875 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 15102 15144 15108 15156
rect 15063 15116 15108 15144
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 17678 15104 17684 15156
rect 17736 15144 17742 15156
rect 19077 15147 19135 15153
rect 19077 15144 19089 15147
rect 17736 15116 19089 15144
rect 17736 15104 17742 15116
rect 19077 15113 19089 15116
rect 19123 15113 19135 15147
rect 19077 15107 19135 15113
rect 20254 15104 20260 15156
rect 20312 15144 20318 15156
rect 20625 15147 20683 15153
rect 20625 15144 20637 15147
rect 20312 15116 20637 15144
rect 20312 15104 20318 15116
rect 20625 15113 20637 15116
rect 20671 15113 20683 15147
rect 20625 15107 20683 15113
rect 20990 15104 20996 15156
rect 21048 15144 21054 15156
rect 22278 15144 22284 15156
rect 21048 15116 22284 15144
rect 21048 15104 21054 15116
rect 22278 15104 22284 15116
rect 22336 15144 22342 15156
rect 23293 15147 23351 15153
rect 22336 15116 23244 15144
rect 22336 15104 22342 15116
rect 12618 15076 12624 15088
rect 12579 15048 12624 15076
rect 12618 15036 12624 15048
rect 12676 15036 12682 15088
rect 13357 15079 13415 15085
rect 13357 15045 13369 15079
rect 13403 15076 13415 15079
rect 13998 15076 14004 15088
rect 13403 15048 14004 15076
rect 13403 15045 13415 15048
rect 13357 15039 13415 15045
rect 13998 15036 14004 15048
rect 14056 15036 14062 15088
rect 17954 15036 17960 15088
rect 18012 15036 18018 15088
rect 18874 15076 18880 15088
rect 18432 15048 18880 15076
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 3421 15011 3479 15017
rect 2832 14980 2877 15008
rect 2832 14968 2838 14980
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 7650 15008 7656 15020
rect 3467 14980 7656 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 15008 12863 15011
rect 13814 15008 13820 15020
rect 12851 14980 13820 15008
rect 12851 14977 12863 14980
rect 12805 14971 12863 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 14977 14427 15011
rect 15194 15008 15200 15020
rect 15155 14980 15200 15008
rect 14369 14971 14427 14977
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 14384 14940 14412 14971
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15562 14968 15568 15020
rect 15620 15008 15626 15020
rect 15657 15011 15715 15017
rect 15657 15008 15669 15011
rect 15620 14980 15669 15008
rect 15620 14968 15626 14980
rect 15657 14977 15669 14980
rect 15703 15008 15715 15011
rect 15703 14980 16528 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 15746 14940 15752 14952
rect 12768 14912 15752 14940
rect 12768 14900 12774 14912
rect 15746 14900 15752 14912
rect 15804 14940 15810 14952
rect 15804 14912 15884 14940
rect 15804 14900 15810 14912
rect 13630 14872 13636 14884
rect 13591 14844 13636 14872
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 15856 14881 15884 14912
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14841 15899 14875
rect 15841 14835 15899 14841
rect 1854 14804 1860 14816
rect 1815 14776 1860 14804
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 3050 14764 3056 14816
rect 3108 14804 3114 14816
rect 3329 14807 3387 14813
rect 3329 14804 3341 14807
rect 3108 14776 3341 14804
rect 3108 14764 3114 14776
rect 3329 14773 3341 14776
rect 3375 14773 3387 14807
rect 14458 14804 14464 14816
rect 14419 14776 14464 14804
rect 3329 14767 3387 14773
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 16500 14804 16528 14980
rect 16666 14940 16672 14952
rect 16627 14912 16672 14940
rect 16666 14900 16672 14912
rect 16724 14900 16730 14952
rect 16945 14943 17003 14949
rect 16945 14909 16957 14943
rect 16991 14940 17003 14943
rect 17310 14940 17316 14952
rect 16991 14912 17316 14940
rect 16991 14909 17003 14912
rect 16945 14903 17003 14909
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18432 14949 18460 15048
rect 18874 15036 18880 15048
rect 18932 15036 18938 15088
rect 20898 15076 20904 15088
rect 20859 15048 20904 15076
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 19426 15008 19432 15020
rect 19260 14980 19432 15008
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 18012 14912 18429 14940
rect 18012 14900 18018 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18417 14903 18475 14909
rect 19260 14881 19288 14980
rect 19426 14968 19432 14980
rect 19484 15008 19490 15020
rect 19705 15011 19763 15017
rect 19705 15008 19717 15011
rect 19484 14980 19717 15008
rect 19484 14968 19490 14980
rect 19705 14977 19717 14980
rect 19751 14977 19763 15011
rect 19886 15008 19892 15020
rect 19847 14980 19892 15008
rect 19705 14971 19763 14977
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 20806 15008 20812 15020
rect 20767 14980 20812 15008
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 20990 15008 20996 15020
rect 20951 14980 20996 15008
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 21111 15011 21169 15017
rect 21111 15008 21123 15011
rect 21109 14977 21123 15008
rect 21157 14977 21169 15011
rect 21109 14971 21169 14977
rect 20070 14900 20076 14952
rect 20128 14940 20134 14952
rect 21109 14940 21137 14971
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 23109 15011 23167 15017
rect 23109 15008 23121 15011
rect 21968 14980 23121 15008
rect 21968 14968 21974 14980
rect 23109 14977 23121 14980
rect 23155 14977 23167 15011
rect 23216 15008 23244 15116
rect 23293 15113 23305 15147
rect 23339 15144 23351 15147
rect 23566 15144 23572 15156
rect 23339 15116 23572 15144
rect 23339 15113 23351 15116
rect 23293 15107 23351 15113
rect 23566 15104 23572 15116
rect 23624 15144 23630 15156
rect 24305 15147 24363 15153
rect 24305 15144 24317 15147
rect 23624 15116 24317 15144
rect 23624 15104 23630 15116
rect 24305 15113 24317 15116
rect 24351 15113 24363 15147
rect 24305 15107 24363 15113
rect 25038 15104 25044 15156
rect 25096 15144 25102 15156
rect 25593 15147 25651 15153
rect 25593 15144 25605 15147
rect 25096 15116 25605 15144
rect 25096 15104 25102 15116
rect 25593 15113 25605 15116
rect 25639 15113 25651 15147
rect 25593 15107 25651 15113
rect 25866 15104 25872 15156
rect 25924 15144 25930 15156
rect 26237 15147 26295 15153
rect 26237 15144 26249 15147
rect 25924 15116 26249 15144
rect 25924 15104 25930 15116
rect 26237 15113 26249 15116
rect 26283 15113 26295 15147
rect 29362 15144 29368 15156
rect 29323 15116 29368 15144
rect 26237 15107 26295 15113
rect 29362 15104 29368 15116
rect 29420 15104 29426 15156
rect 29822 15144 29828 15156
rect 29783 15116 29828 15144
rect 29822 15104 29828 15116
rect 29880 15104 29886 15156
rect 30282 15104 30288 15156
rect 30340 15144 30346 15156
rect 30837 15147 30895 15153
rect 30837 15144 30849 15147
rect 30340 15116 30849 15144
rect 30340 15104 30346 15116
rect 30837 15113 30849 15116
rect 30883 15113 30895 15147
rect 31478 15144 31484 15156
rect 30837 15107 30895 15113
rect 30944 15116 31484 15144
rect 24121 15079 24179 15085
rect 24121 15045 24133 15079
rect 24167 15076 24179 15079
rect 25685 15079 25743 15085
rect 24167 15048 25636 15076
rect 24167 15045 24179 15048
rect 24121 15039 24179 15045
rect 25608 15020 25636 15048
rect 25685 15045 25697 15079
rect 25731 15076 25743 15079
rect 26970 15076 26976 15088
rect 25731 15048 26976 15076
rect 25731 15045 25743 15048
rect 25685 15039 25743 15045
rect 26970 15036 26976 15048
rect 27028 15036 27034 15088
rect 28994 15076 29000 15088
rect 27632 15048 29000 15076
rect 23290 15008 23296 15020
rect 23216 14980 23296 15008
rect 23109 14971 23167 14977
rect 23290 14968 23296 14980
rect 23348 15008 23354 15020
rect 24397 15011 24455 15017
rect 23348 14980 23441 15008
rect 23348 14968 23354 14980
rect 24397 14977 24409 15011
rect 24443 14977 24455 15011
rect 24854 15008 24860 15020
rect 24815 14980 24860 15008
rect 24397 14971 24455 14977
rect 20128 14912 21137 14940
rect 21269 14943 21327 14949
rect 20128 14900 20134 14912
rect 21269 14909 21281 14943
rect 21315 14909 21327 14943
rect 21818 14940 21824 14952
rect 21779 14912 21824 14940
rect 21269 14903 21327 14909
rect 19245 14875 19303 14881
rect 17972 14844 19196 14872
rect 17972 14804 18000 14844
rect 19058 14804 19064 14816
rect 16500 14776 18000 14804
rect 19019 14776 19064 14804
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 19168 14804 19196 14844
rect 19245 14841 19257 14875
rect 19291 14841 19303 14875
rect 19245 14835 19303 14841
rect 19334 14804 19340 14816
rect 19168 14776 19340 14804
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19702 14804 19708 14816
rect 19663 14776 19708 14804
rect 19702 14764 19708 14776
rect 19760 14804 19766 14816
rect 19978 14804 19984 14816
rect 19760 14776 19984 14804
rect 19760 14764 19766 14776
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 21284 14804 21312 14903
rect 21818 14900 21824 14912
rect 21876 14900 21882 14952
rect 22002 14900 22008 14952
rect 22060 14940 22066 14952
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 22060 14912 22109 14940
rect 22060 14900 22066 14912
rect 22097 14909 22109 14912
rect 22143 14909 22155 14943
rect 24412 14940 24440 14971
rect 24854 14968 24860 14980
rect 24912 14968 24918 15020
rect 25041 15011 25099 15017
rect 25041 14977 25053 15011
rect 25087 15008 25099 15011
rect 25087 14980 25544 15008
rect 25087 14977 25099 14980
rect 25041 14971 25099 14977
rect 24949 14943 25007 14949
rect 24949 14940 24961 14943
rect 24412 14912 24961 14940
rect 22097 14903 22155 14909
rect 24949 14909 24961 14912
rect 24995 14909 25007 14943
rect 24949 14903 25007 14909
rect 21726 14832 21732 14884
rect 21784 14872 21790 14884
rect 25222 14872 25228 14884
rect 21784 14844 25228 14872
rect 21784 14832 21790 14844
rect 25222 14832 25228 14844
rect 25280 14832 25286 14884
rect 25314 14832 25320 14884
rect 25372 14872 25378 14884
rect 25516 14872 25544 14980
rect 25590 14968 25596 15020
rect 25648 14968 25654 15020
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26418 15008 26424 15020
rect 26379 14980 26424 15008
rect 26237 14971 26295 14977
rect 26252 14940 26280 14971
rect 26418 14968 26424 14980
rect 26476 14968 26482 15020
rect 27632 15008 27660 15048
rect 28994 15036 29000 15048
rect 29052 15036 29058 15088
rect 30944 15076 30972 15116
rect 31478 15104 31484 15116
rect 31536 15144 31542 15156
rect 32125 15147 32183 15153
rect 32125 15144 32137 15147
rect 31536 15116 32137 15144
rect 31536 15104 31542 15116
rect 32125 15113 32137 15116
rect 32171 15113 32183 15147
rect 32125 15107 32183 15113
rect 32293 15147 32351 15153
rect 32293 15113 32305 15147
rect 32339 15144 32351 15147
rect 32398 15144 32404 15156
rect 32339 15116 32404 15144
rect 32339 15113 32351 15116
rect 32293 15107 32351 15113
rect 32398 15104 32404 15116
rect 32456 15104 32462 15156
rect 36538 15144 36544 15156
rect 33060 15116 36544 15144
rect 31018 15085 31024 15088
rect 29196 15048 30972 15076
rect 31000 15079 31024 15085
rect 26804 14980 27660 15008
rect 27709 15011 27767 15017
rect 26694 14940 26700 14952
rect 26252 14912 26700 14940
rect 26694 14900 26700 14912
rect 26752 14900 26758 14952
rect 26804 14872 26832 14980
rect 27709 14977 27721 15011
rect 27755 15008 27767 15011
rect 27890 15008 27896 15020
rect 27755 14980 27896 15008
rect 27755 14977 27767 14980
rect 27709 14971 27767 14977
rect 27890 14968 27896 14980
rect 27948 14968 27954 15020
rect 29086 15008 29092 15020
rect 28184 14980 29092 15008
rect 27525 14943 27583 14949
rect 27525 14909 27537 14943
rect 27571 14909 27583 14943
rect 27525 14903 27583 14909
rect 27617 14943 27675 14949
rect 27617 14909 27629 14943
rect 27663 14940 27675 14943
rect 27798 14940 27804 14952
rect 27663 14912 27804 14940
rect 27663 14909 27675 14912
rect 27617 14903 27675 14909
rect 25372 14844 26832 14872
rect 27540 14872 27568 14903
rect 27798 14900 27804 14912
rect 27856 14900 27862 14952
rect 28184 14872 28212 14980
rect 29086 14968 29092 14980
rect 29144 14968 29150 15020
rect 29196 15017 29224 15048
rect 31000 15045 31012 15079
rect 31000 15039 31024 15045
rect 31018 15036 31024 15039
rect 31076 15036 31082 15088
rect 31202 15076 31208 15088
rect 31163 15048 31208 15076
rect 31202 15036 31208 15048
rect 31260 15036 31266 15088
rect 32490 15076 32496 15088
rect 32451 15048 32496 15076
rect 32490 15036 32496 15048
rect 32548 15036 32554 15088
rect 29181 15011 29239 15017
rect 29181 14977 29193 15011
rect 29227 14977 29239 15011
rect 29181 14971 29239 14977
rect 29546 14968 29552 15020
rect 29604 15008 29610 15020
rect 30009 15011 30067 15017
rect 30009 15008 30021 15011
rect 29604 14980 30021 15008
rect 29604 14968 29610 14980
rect 30009 14977 30021 14980
rect 30055 14977 30067 15011
rect 30009 14971 30067 14977
rect 30285 15011 30343 15017
rect 30285 14977 30297 15011
rect 30331 15008 30343 15011
rect 30834 15008 30840 15020
rect 30331 14980 30840 15008
rect 30331 14977 30343 14980
rect 30285 14971 30343 14977
rect 30834 14968 30840 14980
rect 30892 14968 30898 15020
rect 31110 14968 31116 15020
rect 31168 15008 31174 15020
rect 31662 15008 31668 15020
rect 31168 14980 31668 15008
rect 31168 14968 31174 14980
rect 31662 14968 31668 14980
rect 31720 15008 31726 15020
rect 33060 15017 33088 15116
rect 36538 15104 36544 15116
rect 36596 15104 36602 15156
rect 33318 15076 33324 15088
rect 33279 15048 33324 15076
rect 33318 15036 33324 15048
rect 33376 15036 33382 15088
rect 34790 15036 34796 15088
rect 34848 15076 34854 15088
rect 35529 15079 35587 15085
rect 35529 15076 35541 15079
rect 34848 15048 35541 15076
rect 34848 15036 34854 15048
rect 35529 15045 35541 15048
rect 35575 15076 35587 15079
rect 35618 15076 35624 15088
rect 35575 15048 35624 15076
rect 35575 15045 35587 15048
rect 35529 15039 35587 15045
rect 35618 15036 35624 15048
rect 35676 15036 35682 15088
rect 36354 15036 36360 15088
rect 36412 15076 36418 15088
rect 36633 15079 36691 15085
rect 36633 15076 36645 15079
rect 36412 15048 36645 15076
rect 36412 15036 36418 15048
rect 36633 15045 36645 15048
rect 36679 15045 36691 15079
rect 36633 15039 36691 15045
rect 33045 15011 33103 15017
rect 33045 15008 33057 15011
rect 31720 14980 33057 15008
rect 31720 14968 31726 14980
rect 33045 14977 33057 14980
rect 33091 14977 33103 15011
rect 33045 14971 33103 14977
rect 34422 14968 34428 15020
rect 34480 14968 34486 15020
rect 35434 15008 35440 15020
rect 35395 14980 35440 15008
rect 35434 14968 35440 14980
rect 35492 14968 35498 15020
rect 35710 15008 35716 15020
rect 35671 14980 35716 15008
rect 35710 14968 35716 14980
rect 35768 14968 35774 15020
rect 35802 14968 35808 15020
rect 35860 15008 35866 15020
rect 36541 15011 36599 15017
rect 36541 15008 36553 15011
rect 35860 14980 36553 15008
rect 35860 14968 35866 14980
rect 36541 14977 36553 14980
rect 36587 14977 36599 15011
rect 36541 14971 36599 14977
rect 37461 15011 37519 15017
rect 37461 14977 37473 15011
rect 37507 15008 37519 15011
rect 38286 15008 38292 15020
rect 37507 14980 38292 15008
rect 37507 14977 37519 14980
rect 37461 14971 37519 14977
rect 38286 14968 38292 14980
rect 38344 14968 38350 15020
rect 28997 14943 29055 14949
rect 28997 14909 29009 14943
rect 29043 14909 29055 14943
rect 28997 14903 29055 14909
rect 30193 14943 30251 14949
rect 30193 14909 30205 14943
rect 30239 14940 30251 14943
rect 31478 14940 31484 14952
rect 30239 14912 31484 14940
rect 30239 14909 30251 14912
rect 30193 14903 30251 14909
rect 27540 14844 28212 14872
rect 29012 14872 29040 14903
rect 31478 14900 31484 14912
rect 31536 14900 31542 14952
rect 32214 14900 32220 14952
rect 32272 14940 32278 14952
rect 34793 14943 34851 14949
rect 34793 14940 34805 14943
rect 32272 14912 34805 14940
rect 32272 14900 32278 14912
rect 34793 14909 34805 14912
rect 34839 14940 34851 14943
rect 35342 14940 35348 14952
rect 34839 14912 35348 14940
rect 34839 14909 34851 14912
rect 34793 14903 34851 14909
rect 35342 14900 35348 14912
rect 35400 14900 35406 14952
rect 29012 14844 30328 14872
rect 25372 14832 25378 14844
rect 21358 14804 21364 14816
rect 21284 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14804 21422 14816
rect 21542 14804 21548 14816
rect 21416 14776 21548 14804
rect 21416 14764 21422 14776
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 24121 14807 24179 14813
rect 24121 14773 24133 14807
rect 24167 14804 24179 14807
rect 25866 14804 25872 14816
rect 24167 14776 25872 14804
rect 24167 14773 24179 14776
rect 24121 14767 24179 14773
rect 25866 14764 25872 14776
rect 25924 14764 25930 14816
rect 28077 14807 28135 14813
rect 28077 14773 28089 14807
rect 28123 14804 28135 14807
rect 28994 14804 29000 14816
rect 28123 14776 29000 14804
rect 28123 14773 28135 14776
rect 28077 14767 28135 14773
rect 28994 14764 29000 14776
rect 29052 14764 29058 14816
rect 30300 14813 30328 14844
rect 35250 14832 35256 14884
rect 35308 14832 35314 14884
rect 30285 14807 30343 14813
rect 30285 14773 30297 14807
rect 30331 14804 30343 14807
rect 30558 14804 30564 14816
rect 30331 14776 30564 14804
rect 30331 14773 30343 14776
rect 30285 14767 30343 14773
rect 30558 14764 30564 14776
rect 30616 14764 30622 14816
rect 31018 14804 31024 14816
rect 30979 14776 31024 14804
rect 31018 14764 31024 14776
rect 31076 14764 31082 14816
rect 32306 14804 32312 14816
rect 32267 14776 32312 14804
rect 32306 14764 32312 14776
rect 32364 14764 32370 14816
rect 32398 14764 32404 14816
rect 32456 14804 32462 14816
rect 33778 14804 33784 14816
rect 32456 14776 33784 14804
rect 32456 14764 32462 14776
rect 33778 14764 33784 14776
rect 33836 14764 33842 14816
rect 35268 14804 35296 14832
rect 35342 14804 35348 14816
rect 35268 14776 35348 14804
rect 35342 14764 35348 14776
rect 35400 14764 35406 14816
rect 35713 14807 35771 14813
rect 35713 14773 35725 14807
rect 35759 14804 35771 14807
rect 35802 14804 35808 14816
rect 35759 14776 35808 14804
rect 35759 14773 35771 14776
rect 35713 14767 35771 14773
rect 35802 14764 35808 14776
rect 35860 14764 35866 14816
rect 36722 14764 36728 14816
rect 36780 14804 36786 14816
rect 37553 14807 37611 14813
rect 37553 14804 37565 14807
rect 36780 14776 37565 14804
rect 36780 14764 36786 14776
rect 37553 14773 37565 14776
rect 37599 14773 37611 14807
rect 37553 14767 37611 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12584 14572 13001 14600
rect 12584 14560 12590 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 17310 14600 17316 14612
rect 17271 14572 17316 14600
rect 12989 14563 13047 14569
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 17494 14560 17500 14612
rect 17552 14600 17558 14612
rect 17681 14603 17739 14609
rect 17681 14600 17693 14603
rect 17552 14572 17693 14600
rect 17552 14560 17558 14572
rect 17681 14569 17693 14572
rect 17727 14569 17739 14603
rect 17681 14563 17739 14569
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 19058 14600 19064 14612
rect 17920 14572 19064 14600
rect 17920 14560 17926 14572
rect 19058 14560 19064 14572
rect 19116 14560 19122 14612
rect 20898 14600 20904 14612
rect 19168 14572 20904 14600
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 14550 14532 14556 14544
rect 2832 14504 14556 14532
rect 2832 14492 2838 14504
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 16853 14535 16911 14541
rect 16853 14501 16865 14535
rect 16899 14532 16911 14535
rect 17218 14532 17224 14544
rect 16899 14504 17224 14532
rect 16899 14501 16911 14504
rect 16853 14495 16911 14501
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 19168 14532 19196 14572
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 21637 14603 21695 14609
rect 21637 14569 21649 14603
rect 21683 14600 21695 14603
rect 21726 14600 21732 14612
rect 21683 14572 21732 14600
rect 21683 14569 21695 14572
rect 21637 14563 21695 14569
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 23290 14560 23296 14612
rect 23348 14600 23354 14612
rect 25406 14600 25412 14612
rect 23348 14572 25412 14600
rect 23348 14560 23354 14572
rect 25406 14560 25412 14572
rect 25464 14560 25470 14612
rect 31665 14603 31723 14609
rect 31665 14569 31677 14603
rect 31711 14600 31723 14603
rect 32306 14600 32312 14612
rect 31711 14572 32312 14600
rect 31711 14569 31723 14572
rect 31665 14563 31723 14569
rect 32306 14560 32312 14572
rect 32364 14560 32370 14612
rect 33781 14603 33839 14609
rect 33781 14569 33793 14603
rect 33827 14600 33839 14603
rect 33870 14600 33876 14612
rect 33827 14572 33876 14600
rect 33827 14569 33839 14572
rect 33781 14563 33839 14569
rect 33870 14560 33876 14572
rect 33928 14560 33934 14612
rect 37458 14600 37464 14612
rect 34532 14572 37464 14600
rect 17328 14504 19196 14532
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 17328 14464 17356 14504
rect 19334 14492 19340 14544
rect 19392 14532 19398 14544
rect 20622 14532 20628 14544
rect 19392 14504 20628 14532
rect 19392 14492 19398 14504
rect 20622 14492 20628 14504
rect 20680 14492 20686 14544
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 21085 14535 21143 14541
rect 21085 14532 21097 14535
rect 20772 14504 21097 14532
rect 20772 14492 20778 14504
rect 21085 14501 21097 14504
rect 21131 14532 21143 14535
rect 21542 14532 21548 14544
rect 21131 14504 21548 14532
rect 21131 14501 21143 14504
rect 21085 14495 21143 14501
rect 21542 14492 21548 14504
rect 21600 14532 21606 14544
rect 24397 14535 24455 14541
rect 24397 14532 24409 14535
rect 21600 14504 24409 14532
rect 21600 14492 21606 14504
rect 24397 14501 24409 14504
rect 24443 14532 24455 14535
rect 24854 14532 24860 14544
rect 24443 14504 24860 14532
rect 24443 14501 24455 14504
rect 24397 14495 24455 14501
rect 24854 14492 24860 14504
rect 24912 14492 24918 14544
rect 30742 14492 30748 14544
rect 30800 14532 30806 14544
rect 30800 14504 31708 14532
rect 30800 14492 30806 14504
rect 19702 14464 19708 14476
rect 15764 14436 17356 14464
rect 17512 14436 19708 14464
rect 15764 14408 15792 14436
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3283 14368 3801 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 13170 14396 13176 14408
rect 13131 14368 13176 14396
rect 3789 14359 3847 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14396 14795 14399
rect 15654 14396 15660 14408
rect 14783 14368 15660 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15746 14356 15752 14408
rect 15804 14396 15810 14408
rect 15804 14368 15897 14396
rect 15804 14356 15810 14368
rect 15930 14356 15936 14408
rect 15988 14396 15994 14408
rect 16577 14399 16635 14405
rect 15988 14368 16033 14396
rect 15988 14356 15994 14368
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 17034 14396 17040 14408
rect 16623 14368 17040 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 17034 14356 17040 14368
rect 17092 14356 17098 14408
rect 17512 14405 17540 14436
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 20533 14467 20591 14473
rect 20533 14433 20545 14467
rect 20579 14464 20591 14467
rect 20806 14464 20812 14476
rect 20579 14436 20812 14464
rect 20579 14433 20591 14436
rect 20533 14427 20591 14433
rect 20806 14424 20812 14436
rect 20864 14464 20870 14476
rect 20864 14436 22508 14464
rect 20864 14424 20870 14436
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 17954 14396 17960 14408
rect 17819 14368 17960 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 18230 14396 18236 14408
rect 18191 14368 18236 14396
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 16853 14331 16911 14337
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 17678 14328 17684 14340
rect 16899 14300 17684 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 17678 14288 17684 14300
rect 17736 14328 17742 14340
rect 18046 14328 18052 14340
rect 17736 14300 18052 14328
rect 17736 14288 17742 14300
rect 18046 14288 18052 14300
rect 18104 14288 18110 14340
rect 18432 14328 18460 14359
rect 18506 14356 18512 14408
rect 18564 14396 18570 14408
rect 18782 14396 18788 14408
rect 18564 14368 18788 14396
rect 18564 14356 18570 14368
rect 18782 14356 18788 14368
rect 18840 14396 18846 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 18840 14368 19625 14396
rect 18840 14356 18846 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 20625 14399 20683 14405
rect 20487 14368 20576 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 18966 14328 18972 14340
rect 18432 14300 18972 14328
rect 18966 14288 18972 14300
rect 19024 14288 19030 14340
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 14240 14232 14657 14260
rect 14240 14220 14246 14232
rect 14645 14229 14657 14232
rect 14691 14229 14703 14263
rect 14645 14223 14703 14229
rect 15933 14263 15991 14269
rect 15933 14229 15945 14263
rect 15979 14260 15991 14263
rect 16574 14260 16580 14272
rect 15979 14232 16580 14260
rect 15979 14229 15991 14232
rect 15933 14223 15991 14229
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 17862 14260 17868 14272
rect 16715 14232 17868 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 18325 14263 18383 14269
rect 18325 14260 18337 14263
rect 18012 14232 18337 14260
rect 18012 14220 18018 14232
rect 18325 14229 18337 14232
rect 18371 14229 18383 14263
rect 18325 14223 18383 14229
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 19521 14263 19579 14269
rect 19521 14260 19533 14263
rect 19484 14232 19533 14260
rect 19484 14220 19490 14232
rect 19521 14229 19533 14232
rect 19567 14229 19579 14263
rect 20548 14260 20576 14368
rect 20625 14365 20637 14399
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14396 21327 14399
rect 21818 14396 21824 14408
rect 21315 14368 21824 14396
rect 21315 14365 21327 14368
rect 21269 14359 21327 14365
rect 20640 14328 20668 14359
rect 21818 14356 21824 14368
rect 21876 14396 21882 14408
rect 22480 14405 22508 14436
rect 22554 14424 22560 14476
rect 22612 14464 22618 14476
rect 23290 14464 23296 14476
rect 22612 14436 22657 14464
rect 22756 14436 23296 14464
rect 22612 14424 22618 14436
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 21876 14368 22201 14396
rect 21876 14356 21882 14368
rect 22189 14365 22201 14368
rect 22235 14396 22247 14399
rect 22465 14399 22523 14405
rect 22235 14368 22324 14396
rect 22235 14365 22247 14368
rect 22189 14359 22247 14365
rect 21726 14328 21732 14340
rect 20640 14300 21404 14328
rect 21376 14272 21404 14300
rect 21468 14300 21732 14328
rect 20990 14260 20996 14272
rect 20548 14232 20996 14260
rect 19521 14223 19579 14229
rect 20990 14220 20996 14232
rect 21048 14220 21054 14272
rect 21358 14260 21364 14272
rect 21319 14232 21364 14260
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 21468 14269 21496 14300
rect 21726 14288 21732 14300
rect 21784 14288 21790 14340
rect 22094 14288 22100 14340
rect 22152 14328 22158 14340
rect 22296 14328 22324 14368
rect 22465 14365 22477 14399
rect 22511 14365 22523 14399
rect 22465 14359 22523 14365
rect 22756 14328 22784 14436
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 23566 14464 23572 14476
rect 23527 14436 23572 14464
rect 23566 14424 23572 14436
rect 23624 14424 23630 14476
rect 25130 14424 25136 14476
rect 25188 14464 25194 14476
rect 26145 14467 26203 14473
rect 26145 14464 26157 14467
rect 25188 14436 26157 14464
rect 25188 14424 25194 14436
rect 26145 14433 26157 14436
rect 26191 14464 26203 14467
rect 27065 14467 27123 14473
rect 27065 14464 27077 14467
rect 26191 14436 27077 14464
rect 26191 14433 26203 14436
rect 26145 14427 26203 14433
rect 27065 14433 27077 14436
rect 27111 14433 27123 14467
rect 27065 14427 27123 14433
rect 28813 14467 28871 14473
rect 28813 14433 28825 14467
rect 28859 14464 28871 14467
rect 29546 14464 29552 14476
rect 28859 14436 29552 14464
rect 28859 14433 28871 14436
rect 28813 14427 28871 14433
rect 29546 14424 29552 14436
rect 29604 14424 29610 14476
rect 29825 14467 29883 14473
rect 29825 14433 29837 14467
rect 29871 14464 29883 14467
rect 30282 14464 30288 14476
rect 29871 14436 30288 14464
rect 29871 14433 29883 14436
rect 29825 14427 29883 14433
rect 30282 14424 30288 14436
rect 30340 14424 30346 14476
rect 31113 14467 31171 14473
rect 31113 14433 31125 14467
rect 31159 14464 31171 14467
rect 31478 14464 31484 14476
rect 31159 14436 31484 14464
rect 31159 14433 31171 14436
rect 31113 14427 31171 14433
rect 31478 14424 31484 14436
rect 31536 14424 31542 14476
rect 31680 14464 31708 14504
rect 31754 14492 31760 14544
rect 31812 14532 31818 14544
rect 34532 14532 34560 14572
rect 37458 14560 37464 14572
rect 37516 14560 37522 14612
rect 31812 14504 34560 14532
rect 31812 14492 31818 14504
rect 34606 14492 34612 14544
rect 34664 14532 34670 14544
rect 35342 14532 35348 14544
rect 34664 14504 35348 14532
rect 34664 14492 34670 14504
rect 35342 14492 35348 14504
rect 35400 14492 35406 14544
rect 32401 14467 32459 14473
rect 32401 14464 32413 14467
rect 31680 14436 32413 14464
rect 32401 14433 32413 14436
rect 32447 14433 32459 14467
rect 32401 14427 32459 14433
rect 36449 14467 36507 14473
rect 36449 14433 36461 14467
rect 36495 14464 36507 14467
rect 36722 14464 36728 14476
rect 36495 14436 36728 14464
rect 36495 14433 36507 14436
rect 36449 14427 36507 14433
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 22152 14300 22197 14328
rect 22296 14300 22784 14328
rect 23032 14368 23397 14396
rect 22152 14288 22158 14300
rect 21453 14263 21511 14269
rect 21453 14229 21465 14263
rect 21499 14229 21511 14263
rect 21453 14223 21511 14229
rect 22741 14263 22799 14269
rect 22741 14229 22753 14263
rect 22787 14260 22799 14263
rect 23032 14260 23060 14368
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 30834 14356 30840 14408
rect 30892 14396 30898 14408
rect 31202 14396 31208 14408
rect 30892 14368 31208 14396
rect 30892 14356 30898 14368
rect 31202 14356 31208 14368
rect 31260 14396 31266 14408
rect 31297 14399 31355 14405
rect 31297 14396 31309 14399
rect 31260 14368 31309 14396
rect 31260 14356 31266 14368
rect 31297 14365 31309 14368
rect 31343 14365 31355 14399
rect 31297 14359 31355 14365
rect 32030 14356 32036 14408
rect 32088 14396 32094 14408
rect 32125 14399 32183 14405
rect 32125 14396 32137 14399
rect 32088 14368 32137 14396
rect 32088 14356 32094 14368
rect 32125 14365 32137 14368
rect 32171 14365 32183 14399
rect 32416 14396 32444 14427
rect 36722 14424 36728 14436
rect 36780 14424 36786 14476
rect 38102 14464 38108 14476
rect 38063 14436 38108 14464
rect 38102 14424 38108 14436
rect 38160 14424 38166 14476
rect 34146 14396 34152 14408
rect 32416 14368 34152 14396
rect 32125 14359 32183 14365
rect 33735 14365 33793 14368
rect 23658 14288 23664 14340
rect 23716 14328 23722 14340
rect 25866 14328 25872 14340
rect 23716 14300 24702 14328
rect 25827 14300 25872 14328
rect 23716 14288 23722 14300
rect 25866 14288 25872 14300
rect 25924 14288 25930 14340
rect 27341 14331 27399 14337
rect 27341 14297 27353 14331
rect 27387 14297 27399 14331
rect 27341 14291 27399 14297
rect 22787 14232 23060 14260
rect 23201 14263 23259 14269
rect 22787 14229 22799 14232
rect 22741 14223 22799 14229
rect 23201 14229 23213 14263
rect 23247 14260 23259 14263
rect 23382 14260 23388 14272
rect 23247 14232 23388 14260
rect 23247 14229 23259 14232
rect 23201 14223 23259 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 27356 14260 27384 14291
rect 27430 14288 27436 14340
rect 27488 14328 27494 14340
rect 31481 14331 31539 14337
rect 27488 14300 27830 14328
rect 27488 14288 27494 14300
rect 31481 14297 31493 14331
rect 31527 14328 31539 14331
rect 32214 14328 32220 14340
rect 31527 14300 32220 14328
rect 31527 14297 31539 14300
rect 31481 14291 31539 14297
rect 32214 14288 32220 14300
rect 32272 14288 32278 14340
rect 33735 14331 33747 14365
rect 33781 14331 33793 14365
rect 34146 14356 34152 14368
rect 34204 14356 34210 14408
rect 36170 14356 36176 14408
rect 36228 14396 36234 14408
rect 36265 14399 36323 14405
rect 36265 14396 36277 14399
rect 36228 14368 36277 14396
rect 36228 14356 36234 14368
rect 36265 14365 36277 14368
rect 36311 14365 36323 14399
rect 36265 14359 36323 14365
rect 33735 14325 33793 14331
rect 33962 14288 33968 14340
rect 34020 14328 34026 14340
rect 35158 14328 35164 14340
rect 34020 14300 34065 14328
rect 35119 14300 35164 14328
rect 34020 14288 34026 14300
rect 35158 14288 35164 14300
rect 35216 14288 35222 14340
rect 28810 14260 28816 14272
rect 27356 14232 28816 14260
rect 28810 14220 28816 14232
rect 28868 14220 28874 14272
rect 31389 14263 31447 14269
rect 31389 14229 31401 14263
rect 31435 14260 31447 14263
rect 31570 14260 31576 14272
rect 31435 14232 31576 14260
rect 31435 14229 31447 14232
rect 31389 14223 31447 14229
rect 31570 14220 31576 14232
rect 31628 14220 31634 14272
rect 33594 14260 33600 14272
rect 33555 14232 33600 14260
rect 33594 14220 33600 14232
rect 33652 14220 33658 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 12621 14059 12679 14065
rect 12621 14025 12633 14059
rect 12667 14056 12679 14059
rect 13998 14056 14004 14068
rect 12667 14028 14004 14056
rect 12667 14025 12679 14028
rect 12621 14019 12679 14025
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 17589 14059 17647 14065
rect 17589 14056 17601 14059
rect 15252 14028 17601 14056
rect 15252 14016 15258 14028
rect 17589 14025 17601 14028
rect 17635 14025 17647 14059
rect 19334 14056 19340 14068
rect 17589 14019 17647 14025
rect 17696 14028 19340 14056
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 14274 13988 14280 14000
rect 13403 13960 14280 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14458 13948 14464 14000
rect 14516 13988 14522 14000
rect 17218 13988 17224 14000
rect 14516 13960 14674 13988
rect 17179 13960 17224 13988
rect 14516 13948 14522 13960
rect 17218 13948 17224 13960
rect 17276 13948 17282 14000
rect 17405 13991 17463 13997
rect 17405 13957 17417 13991
rect 17451 13988 17463 13991
rect 17494 13988 17500 14000
rect 17451 13960 17500 13988
rect 17451 13957 17463 13960
rect 17405 13951 17463 13957
rect 17494 13948 17500 13960
rect 17552 13948 17558 14000
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 12710 13920 12716 13932
rect 12671 13892 12716 13920
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 13906 13920 13912 13932
rect 13867 13892 13912 13920
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 17696 13920 17724 14028
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 21910 14016 21916 14068
rect 21968 14056 21974 14068
rect 22189 14059 22247 14065
rect 22189 14056 22201 14059
rect 21968 14028 22201 14056
rect 21968 14016 21974 14028
rect 22189 14025 22201 14028
rect 22235 14025 22247 14059
rect 25038 14056 25044 14068
rect 22189 14019 22247 14025
rect 22940 14028 25044 14056
rect 20806 13988 20812 14000
rect 18524 13960 20812 13988
rect 18414 13920 18420 13932
rect 15396 13892 17724 13920
rect 18375 13892 18420 13920
rect 2038 13852 2044 13864
rect 1999 13824 2044 13852
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 13173 13855 13231 13861
rect 2832 13824 2877 13852
rect 2832 13812 2838 13824
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13814 13852 13820 13864
rect 13219 13824 13820 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 14182 13852 14188 13864
rect 14143 13824 14188 13852
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 15396 13852 15424 13892
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 18524 13929 18552 13960
rect 20806 13948 20812 13960
rect 20864 13948 20870 14000
rect 21818 13988 21824 14000
rect 21652 13960 21824 13988
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13889 18567 13923
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 18509 13883 18567 13889
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20162 13920 20168 13932
rect 19935 13892 20168 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20162 13880 20168 13892
rect 20220 13920 20226 13932
rect 20438 13920 20444 13932
rect 20220 13892 20444 13920
rect 20220 13880 20226 13892
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 14608 13824 15424 13852
rect 15657 13855 15715 13861
rect 14608 13812 14614 13824
rect 15657 13821 15669 13855
rect 15703 13852 15715 13855
rect 15930 13852 15936 13864
rect 15703 13824 15936 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 16758 13812 16764 13864
rect 16816 13852 16822 13864
rect 18233 13855 18291 13861
rect 18233 13852 18245 13855
rect 16816 13824 18245 13852
rect 16816 13812 16822 13824
rect 18233 13821 18245 13824
rect 18279 13821 18291 13855
rect 18598 13852 18604 13864
rect 18559 13824 18604 13852
rect 18233 13815 18291 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 19058 13812 19064 13864
rect 19116 13852 19122 13864
rect 20640 13852 20668 13883
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20901 13923 20959 13929
rect 20772 13892 20817 13920
rect 20772 13880 20778 13892
rect 20901 13889 20913 13923
rect 20947 13920 20959 13923
rect 21652 13920 21680 13960
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 22051 13957 22109 13963
rect 22051 13932 22063 13957
rect 20947 13892 21680 13920
rect 20947 13889 20959 13892
rect 20901 13883 20959 13889
rect 21726 13880 21732 13932
rect 21784 13920 21790 13932
rect 22002 13920 22008 13932
rect 21784 13892 22008 13920
rect 21784 13880 21790 13892
rect 22002 13880 22008 13892
rect 22060 13923 22063 13932
rect 22097 13923 22109 13957
rect 22940 13929 22968 14028
rect 25038 14016 25044 14028
rect 25096 14016 25102 14068
rect 25314 14056 25320 14068
rect 25275 14028 25320 14056
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 27801 14059 27859 14065
rect 27801 14025 27813 14059
rect 27847 14056 27859 14059
rect 27890 14056 27896 14068
rect 27847 14028 27896 14056
rect 27847 14025 27859 14028
rect 27801 14019 27859 14025
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 28445 14059 28503 14065
rect 28445 14025 28457 14059
rect 28491 14056 28503 14059
rect 29546 14056 29552 14068
rect 28491 14028 29552 14056
rect 28491 14025 28503 14028
rect 28445 14019 28503 14025
rect 29546 14016 29552 14028
rect 29604 14056 29610 14068
rect 30558 14056 30564 14068
rect 29604 14028 30564 14056
rect 29604 14016 29610 14028
rect 30558 14016 30564 14028
rect 30616 14016 30622 14068
rect 31018 14056 31024 14068
rect 30979 14028 31024 14056
rect 31018 14016 31024 14028
rect 31076 14016 31082 14068
rect 31202 14016 31208 14068
rect 31260 14056 31266 14068
rect 31389 14059 31447 14065
rect 31389 14056 31401 14059
rect 31260 14028 31401 14056
rect 31260 14016 31266 14028
rect 31389 14025 31401 14028
rect 31435 14025 31447 14059
rect 31389 14019 31447 14025
rect 34977 14059 35035 14065
rect 34977 14025 34989 14059
rect 35023 14056 35035 14059
rect 35710 14056 35716 14068
rect 35023 14028 35716 14056
rect 35023 14025 35035 14028
rect 34977 14019 35035 14025
rect 35710 14016 35716 14028
rect 35768 14016 35774 14068
rect 37553 14059 37611 14065
rect 37553 14025 37565 14059
rect 37599 14056 37611 14059
rect 37918 14056 37924 14068
rect 37599 14028 37924 14056
rect 37599 14025 37611 14028
rect 37553 14019 37611 14025
rect 37918 14016 37924 14028
rect 37976 14016 37982 14068
rect 26694 13988 26700 14000
rect 24426 13960 26700 13988
rect 26694 13948 26700 13960
rect 26752 13948 26758 14000
rect 27338 13948 27344 14000
rect 27396 13988 27402 14000
rect 27433 13991 27491 13997
rect 27433 13988 27445 13991
rect 27396 13960 27445 13988
rect 27396 13948 27402 13960
rect 27433 13957 27445 13960
rect 27479 13957 27491 13991
rect 27433 13951 27491 13957
rect 27649 13991 27707 13997
rect 27649 13957 27661 13991
rect 27695 13988 27707 13991
rect 28626 13988 28632 14000
rect 27695 13960 28632 13988
rect 27695 13957 27707 13960
rect 27649 13951 27707 13957
rect 28626 13948 28632 13960
rect 28684 13948 28690 14000
rect 31110 13988 31116 14000
rect 30208 13960 31116 13988
rect 22060 13917 22109 13923
rect 22925 13923 22983 13929
rect 22060 13892 22094 13917
rect 22060 13880 22066 13892
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 25498 13920 25504 13932
rect 25459 13892 25504 13920
rect 22925 13883 22983 13889
rect 25498 13880 25504 13892
rect 25556 13880 25562 13932
rect 26142 13920 26148 13932
rect 26103 13892 26148 13920
rect 26142 13880 26148 13892
rect 26200 13880 26206 13932
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 30208 13929 30236 13960
rect 31110 13948 31116 13960
rect 31168 13948 31174 14000
rect 31570 13988 31576 14000
rect 31312 13960 31576 13988
rect 30193 13923 30251 13929
rect 26292 13892 28842 13920
rect 26292 13880 26298 13892
rect 30193 13889 30205 13923
rect 30239 13889 30251 13923
rect 31202 13920 31208 13932
rect 31163 13892 31208 13920
rect 30193 13883 30251 13889
rect 31202 13880 31208 13892
rect 31260 13880 31266 13932
rect 31312 13929 31340 13960
rect 31570 13948 31576 13960
rect 31628 13948 31634 14000
rect 33152 13960 34100 13988
rect 31297 13923 31355 13929
rect 31297 13889 31309 13923
rect 31343 13889 31355 13923
rect 31297 13883 31355 13889
rect 19116 13824 20668 13852
rect 19116 13812 19122 13824
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 23198 13852 23204 13864
rect 20864 13824 23060 13852
rect 23159 13824 23204 13852
rect 20864 13812 20870 13824
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 10410 13784 10416 13796
rect 5132 13756 10416 13784
rect 5132 13744 5138 13756
rect 10410 13744 10416 13756
rect 10468 13744 10474 13796
rect 15948 13784 15976 13812
rect 17310 13784 17316 13796
rect 15948 13756 17316 13784
rect 17310 13744 17316 13756
rect 17368 13744 17374 13796
rect 19334 13744 19340 13796
rect 19392 13784 19398 13796
rect 19705 13787 19763 13793
rect 19705 13784 19717 13787
rect 19392 13756 19717 13784
rect 19392 13744 19398 13756
rect 19705 13753 19717 13756
rect 19751 13784 19763 13787
rect 19978 13784 19984 13796
rect 19751 13756 19984 13784
rect 19751 13753 19763 13756
rect 19705 13747 19763 13753
rect 19978 13744 19984 13756
rect 20036 13784 20042 13796
rect 21818 13784 21824 13796
rect 20036 13756 21824 13784
rect 20036 13744 20042 13756
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 19242 13716 19248 13728
rect 15528 13688 19248 13716
rect 15528 13676 15534 13688
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 20438 13716 20444 13728
rect 20399 13688 20444 13716
rect 20438 13676 20444 13688
rect 20496 13676 20502 13728
rect 20622 13716 20628 13728
rect 20583 13688 20628 13716
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 22005 13719 22063 13725
rect 22005 13716 22017 13719
rect 21416 13688 22017 13716
rect 21416 13676 21422 13688
rect 22005 13685 22017 13688
rect 22051 13685 22063 13719
rect 23032 13716 23060 13824
rect 23198 13812 23204 13824
rect 23256 13812 23262 13864
rect 23290 13812 23296 13864
rect 23348 13852 23354 13864
rect 24673 13855 24731 13861
rect 24673 13852 24685 13855
rect 23348 13824 24685 13852
rect 23348 13812 23354 13824
rect 24673 13821 24685 13824
rect 24719 13821 24731 13855
rect 24673 13815 24731 13821
rect 28626 13812 28632 13864
rect 28684 13852 28690 13864
rect 29362 13852 29368 13864
rect 28684 13824 29368 13852
rect 28684 13812 28690 13824
rect 29362 13812 29368 13824
rect 29420 13812 29426 13864
rect 29914 13852 29920 13864
rect 29875 13824 29920 13852
rect 29914 13812 29920 13824
rect 29972 13812 29978 13864
rect 31110 13812 31116 13864
rect 31168 13852 31174 13864
rect 31312 13852 31340 13883
rect 32030 13880 32036 13932
rect 32088 13920 32094 13932
rect 32493 13923 32551 13929
rect 32493 13920 32505 13923
rect 32088 13892 32505 13920
rect 32088 13880 32094 13892
rect 32493 13889 32505 13892
rect 32539 13889 32551 13923
rect 32493 13883 32551 13889
rect 32769 13923 32827 13929
rect 32769 13889 32781 13923
rect 32815 13920 32827 13923
rect 32950 13920 32956 13932
rect 32815 13892 32956 13920
rect 32815 13889 32827 13892
rect 32769 13883 32827 13889
rect 32950 13880 32956 13892
rect 33008 13880 33014 13932
rect 31570 13852 31576 13864
rect 31168 13824 31340 13852
rect 31531 13824 31576 13852
rect 31168 13812 31174 13824
rect 31570 13812 31576 13824
rect 31628 13812 31634 13864
rect 33152 13784 33180 13960
rect 33226 13880 33232 13932
rect 33284 13920 33290 13932
rect 34072 13929 34100 13960
rect 35434 13948 35440 14000
rect 35492 13948 35498 14000
rect 36538 13948 36544 14000
rect 36596 13988 36602 14000
rect 36596 13960 36768 13988
rect 36596 13948 36602 13960
rect 33781 13923 33839 13929
rect 33781 13920 33793 13923
rect 33284 13892 33793 13920
rect 33284 13880 33290 13892
rect 33781 13889 33793 13892
rect 33827 13889 33839 13923
rect 33781 13883 33839 13889
rect 34057 13923 34115 13929
rect 34057 13889 34069 13923
rect 34103 13889 34115 13923
rect 34057 13883 34115 13889
rect 34146 13880 34152 13932
rect 34204 13920 34210 13932
rect 36740 13929 36768 13960
rect 36725 13923 36783 13929
rect 34204 13892 34249 13920
rect 34204 13880 34210 13892
rect 36725 13889 36737 13923
rect 36771 13889 36783 13923
rect 37458 13920 37464 13932
rect 37419 13892 37464 13920
rect 36725 13883 36783 13889
rect 37458 13880 37464 13892
rect 37516 13880 37522 13932
rect 33870 13852 33876 13864
rect 33831 13824 33876 13852
rect 33870 13812 33876 13824
rect 33928 13812 33934 13864
rect 34333 13855 34391 13861
rect 34333 13821 34345 13855
rect 34379 13852 34391 13855
rect 35710 13852 35716 13864
rect 34379 13824 35716 13852
rect 34379 13821 34391 13824
rect 34333 13815 34391 13821
rect 35710 13812 35716 13824
rect 35768 13812 35774 13864
rect 36446 13852 36452 13864
rect 36407 13824 36452 13852
rect 36446 13812 36452 13824
rect 36504 13812 36510 13864
rect 32600 13756 33180 13784
rect 32600 13728 32628 13756
rect 24762 13716 24768 13728
rect 23032 13688 24768 13716
rect 22005 13679 22063 13685
rect 24762 13676 24768 13688
rect 24820 13716 24826 13728
rect 26329 13719 26387 13725
rect 26329 13716 26341 13719
rect 24820 13688 26341 13716
rect 24820 13676 24826 13688
rect 26329 13685 26341 13688
rect 26375 13716 26387 13719
rect 27154 13716 27160 13728
rect 26375 13688 27160 13716
rect 26375 13685 26387 13688
rect 26329 13679 26387 13685
rect 27154 13676 27160 13688
rect 27212 13676 27218 13728
rect 27617 13719 27675 13725
rect 27617 13685 27629 13719
rect 27663 13716 27675 13719
rect 27982 13716 27988 13728
rect 27663 13688 27988 13716
rect 27663 13685 27675 13688
rect 27617 13679 27675 13685
rect 27982 13676 27988 13688
rect 28040 13676 28046 13728
rect 29546 13676 29552 13728
rect 29604 13716 29610 13728
rect 32582 13716 32588 13728
rect 29604 13688 32588 13716
rect 29604 13676 29610 13688
rect 32582 13676 32588 13688
rect 32640 13676 32646 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 2501 13515 2559 13521
rect 2501 13512 2513 13515
rect 2096 13484 2513 13512
rect 2096 13472 2102 13484
rect 2501 13481 2513 13484
rect 2547 13481 2559 13515
rect 2501 13475 2559 13481
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 15470 13512 15476 13524
rect 4120 13484 15476 13512
rect 4120 13472 4126 13484
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 15654 13472 15660 13524
rect 15712 13512 15718 13524
rect 16853 13515 16911 13521
rect 16853 13512 16865 13515
rect 15712 13484 16865 13512
rect 15712 13472 15718 13484
rect 16853 13481 16865 13484
rect 16899 13481 16911 13515
rect 18046 13512 18052 13524
rect 18007 13484 18052 13512
rect 16853 13475 16911 13481
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 20346 13512 20352 13524
rect 20307 13484 20352 13512
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21729 13515 21787 13521
rect 21729 13512 21741 13515
rect 21140 13484 21741 13512
rect 21140 13472 21146 13484
rect 21729 13481 21741 13484
rect 21775 13481 21787 13515
rect 23198 13512 23204 13524
rect 23159 13484 23204 13512
rect 21729 13475 21787 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 24949 13515 25007 13521
rect 24949 13481 24961 13515
rect 24995 13512 25007 13515
rect 26234 13512 26240 13524
rect 24995 13484 26240 13512
rect 24995 13481 25007 13484
rect 24949 13475 25007 13481
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 27801 13515 27859 13521
rect 27801 13481 27813 13515
rect 27847 13512 27859 13515
rect 27890 13512 27896 13524
rect 27847 13484 27896 13512
rect 27847 13481 27859 13484
rect 27801 13475 27859 13481
rect 27890 13472 27896 13484
rect 27948 13512 27954 13524
rect 28534 13512 28540 13524
rect 27948 13484 28540 13512
rect 27948 13472 27954 13484
rect 28534 13472 28540 13484
rect 28592 13472 28598 13524
rect 29638 13512 29644 13524
rect 29551 13484 29644 13512
rect 29638 13472 29644 13484
rect 29696 13512 29702 13524
rect 29696 13484 29868 13512
rect 29696 13472 29702 13484
rect 20622 13444 20628 13456
rect 18616 13416 20628 13444
rect 16393 13379 16451 13385
rect 16393 13345 16405 13379
rect 16439 13376 16451 13379
rect 16666 13376 16672 13388
rect 16439 13348 16672 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 17310 13376 17316 13388
rect 17271 13348 17316 13376
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 17494 13376 17500 13388
rect 17455 13348 17500 13376
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 1452 13280 1593 13308
rect 1452 13268 1458 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13308 2651 13311
rect 5074 13308 5080 13320
rect 2639 13280 5080 13308
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 16632 13280 17233 13308
rect 16632 13268 16638 13280
rect 17221 13277 17233 13280
rect 17267 13277 17279 13311
rect 17328 13308 17356 13336
rect 18616 13317 18644 13416
rect 20622 13404 20628 13416
rect 20680 13404 20686 13456
rect 21913 13447 21971 13453
rect 21913 13413 21925 13447
rect 21959 13444 21971 13447
rect 25590 13444 25596 13456
rect 21959 13416 25596 13444
rect 21959 13413 21971 13416
rect 21913 13407 21971 13413
rect 25590 13404 25596 13416
rect 25648 13404 25654 13456
rect 26510 13404 26516 13456
rect 26568 13444 26574 13456
rect 26878 13444 26884 13456
rect 26568 13416 26884 13444
rect 26568 13404 26574 13416
rect 26878 13404 26884 13416
rect 26936 13444 26942 13456
rect 26936 13416 27660 13444
rect 26936 13404 26942 13416
rect 20990 13376 20996 13388
rect 20903 13348 20996 13376
rect 20990 13336 20996 13348
rect 21048 13376 21054 13388
rect 21726 13376 21732 13388
rect 21048 13348 21732 13376
rect 21048 13336 21054 13348
rect 21726 13336 21732 13348
rect 21784 13336 21790 13388
rect 21818 13336 21824 13388
rect 21876 13376 21882 13388
rect 27632 13376 27660 13416
rect 29270 13376 29276 13388
rect 21876 13348 27184 13376
rect 21876 13336 21882 13348
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 17328 13280 18613 13308
rect 17221 13271 17279 13277
rect 18601 13277 18613 13280
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 20346 13308 20352 13320
rect 19659 13280 20352 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 20346 13268 20352 13280
rect 20404 13308 20410 13320
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 20404 13280 20821 13308
rect 20404 13268 20410 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 22370 13268 22376 13320
rect 22428 13308 22434 13320
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 22428 13280 22477 13308
rect 22428 13268 22434 13280
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 22554 13268 22560 13320
rect 22612 13308 22618 13320
rect 22649 13311 22707 13317
rect 22649 13308 22661 13311
rect 22612 13280 22661 13308
rect 22612 13268 22618 13280
rect 22649 13277 22661 13280
rect 22695 13277 22707 13311
rect 23382 13308 23388 13320
rect 23343 13280 23388 13308
rect 22649 13271 22707 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13308 24915 13311
rect 24946 13308 24952 13320
rect 24903 13280 24952 13308
rect 24903 13277 24915 13280
rect 24857 13271 24915 13277
rect 24946 13268 24952 13280
rect 25004 13308 25010 13320
rect 25004 13280 25728 13308
rect 25004 13268 25010 13280
rect 13998 13200 14004 13252
rect 14056 13240 14062 13252
rect 16114 13240 16120 13252
rect 14056 13212 14950 13240
rect 16075 13212 16120 13240
rect 14056 13200 14062 13212
rect 16114 13200 16120 13212
rect 16172 13200 16178 13252
rect 18230 13240 18236 13252
rect 18191 13212 18236 13240
rect 18230 13200 18236 13212
rect 18288 13200 18294 13252
rect 18417 13243 18475 13249
rect 18417 13209 18429 13243
rect 18463 13240 18475 13243
rect 20990 13240 20996 13252
rect 18463 13212 20996 13240
rect 18463 13209 18475 13212
rect 18417 13203 18475 13209
rect 20990 13200 20996 13212
rect 21048 13200 21054 13252
rect 21542 13240 21548 13252
rect 21503 13212 21548 13240
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 21761 13243 21819 13249
rect 21761 13209 21773 13243
rect 21807 13240 21819 13243
rect 21910 13240 21916 13252
rect 21807 13212 21916 13240
rect 21807 13209 21819 13212
rect 21761 13203 21819 13209
rect 21910 13200 21916 13212
rect 21968 13200 21974 13252
rect 22094 13200 22100 13252
rect 22152 13240 22158 13252
rect 23014 13240 23020 13252
rect 22152 13212 23020 13240
rect 22152 13200 22158 13212
rect 23014 13200 23020 13212
rect 23072 13240 23078 13252
rect 23290 13240 23296 13252
rect 23072 13212 23296 13240
rect 23072 13200 23078 13212
rect 23290 13200 23296 13212
rect 23348 13200 23354 13252
rect 23474 13200 23480 13252
rect 23532 13240 23538 13252
rect 25498 13240 25504 13252
rect 23532 13212 25504 13240
rect 23532 13200 23538 13212
rect 25498 13200 25504 13212
rect 25556 13240 25562 13252
rect 25593 13243 25651 13249
rect 25593 13240 25605 13243
rect 25556 13212 25605 13240
rect 25556 13200 25562 13212
rect 25593 13209 25605 13212
rect 25639 13209 25651 13243
rect 25700 13240 25728 13280
rect 25774 13268 25780 13320
rect 25832 13308 25838 13320
rect 26436 13317 26464 13348
rect 26237 13311 26295 13317
rect 26237 13308 26249 13311
rect 25832 13280 26249 13308
rect 25832 13268 25838 13280
rect 26237 13277 26249 13280
rect 26283 13277 26295 13311
rect 26237 13271 26295 13277
rect 26421 13311 26479 13317
rect 26421 13277 26433 13311
rect 26467 13277 26479 13311
rect 26878 13308 26884 13320
rect 26839 13280 26884 13308
rect 26421 13271 26479 13277
rect 26878 13268 26884 13280
rect 26936 13268 26942 13320
rect 25700 13212 27108 13240
rect 25593 13203 25651 13209
rect 27080 13184 27108 13212
rect 14645 13175 14703 13181
rect 14645 13141 14657 13175
rect 14691 13172 14703 13175
rect 16758 13172 16764 13184
rect 14691 13144 16764 13172
rect 14691 13141 14703 13144
rect 14645 13135 14703 13141
rect 16758 13132 16764 13144
rect 16816 13132 16822 13184
rect 18322 13172 18328 13184
rect 18283 13144 18328 13172
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 19797 13175 19855 13181
rect 19797 13141 19809 13175
rect 19843 13172 19855 13175
rect 19978 13172 19984 13184
rect 19843 13144 19984 13172
rect 19843 13141 19855 13144
rect 19797 13135 19855 13141
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 22462 13172 22468 13184
rect 22244 13144 22468 13172
rect 22244 13132 22250 13144
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 22649 13175 22707 13181
rect 22649 13141 22661 13175
rect 22695 13172 22707 13175
rect 24302 13172 24308 13184
rect 22695 13144 24308 13172
rect 22695 13141 22707 13144
rect 22649 13135 22707 13141
rect 24302 13132 24308 13144
rect 24360 13172 24366 13184
rect 24762 13172 24768 13184
rect 24360 13144 24768 13172
rect 24360 13132 24366 13144
rect 24762 13132 24768 13144
rect 24820 13132 24826 13184
rect 25682 13172 25688 13184
rect 25643 13144 25688 13172
rect 25682 13132 25688 13144
rect 25740 13172 25746 13184
rect 26050 13172 26056 13184
rect 25740 13144 26056 13172
rect 25740 13132 25746 13144
rect 26050 13132 26056 13144
rect 26108 13132 26114 13184
rect 26326 13172 26332 13184
rect 26287 13144 26332 13172
rect 26326 13132 26332 13144
rect 26384 13132 26390 13184
rect 27062 13172 27068 13184
rect 27023 13144 27068 13172
rect 27062 13132 27068 13144
rect 27120 13132 27126 13184
rect 27156 13172 27184 13348
rect 27632 13348 29276 13376
rect 27632 13317 27660 13348
rect 29270 13336 29276 13348
rect 29328 13336 29334 13388
rect 29454 13336 29460 13388
rect 29512 13376 29518 13388
rect 29549 13379 29607 13385
rect 29549 13376 29561 13379
rect 29512 13348 29561 13376
rect 29512 13336 29518 13348
rect 29549 13345 29561 13348
rect 29595 13345 29607 13379
rect 29840 13376 29868 13484
rect 29914 13472 29920 13524
rect 29972 13512 29978 13524
rect 30009 13515 30067 13521
rect 30009 13512 30021 13515
rect 29972 13484 30021 13512
rect 29972 13472 29978 13484
rect 30009 13481 30021 13484
rect 30055 13481 30067 13515
rect 30009 13475 30067 13481
rect 30650 13472 30656 13524
rect 30708 13512 30714 13524
rect 33689 13515 33747 13521
rect 33689 13512 33701 13515
rect 30708 13484 33701 13512
rect 30708 13472 30714 13484
rect 33689 13481 33701 13484
rect 33735 13481 33747 13515
rect 34146 13512 34152 13524
rect 34107 13484 34152 13512
rect 33689 13475 33747 13481
rect 34146 13472 34152 13484
rect 34204 13472 34210 13524
rect 33870 13404 33876 13456
rect 33928 13444 33934 13456
rect 34054 13444 34060 13456
rect 33928 13416 34060 13444
rect 33928 13404 33934 13416
rect 34054 13404 34060 13416
rect 34112 13444 34118 13456
rect 34701 13447 34759 13453
rect 34701 13444 34713 13447
rect 34112 13416 34713 13444
rect 34112 13404 34118 13416
rect 34701 13413 34713 13416
rect 34747 13444 34759 13447
rect 35158 13444 35164 13456
rect 34747 13416 35164 13444
rect 34747 13413 34759 13416
rect 34701 13407 34759 13413
rect 35158 13404 35164 13416
rect 35216 13404 35222 13456
rect 30929 13379 30987 13385
rect 30929 13376 30941 13379
rect 29840 13348 30941 13376
rect 29549 13339 29607 13345
rect 30929 13345 30941 13348
rect 30975 13345 30987 13379
rect 30929 13339 30987 13345
rect 31018 13336 31024 13388
rect 31076 13376 31082 13388
rect 31297 13379 31355 13385
rect 31297 13376 31309 13379
rect 31076 13348 31309 13376
rect 31076 13336 31082 13348
rect 31297 13345 31309 13348
rect 31343 13345 31355 13379
rect 31297 13339 31355 13345
rect 32490 13336 32496 13388
rect 32548 13376 32554 13388
rect 32861 13379 32919 13385
rect 32861 13376 32873 13379
rect 32548 13348 32873 13376
rect 32548 13336 32554 13348
rect 32861 13345 32873 13348
rect 32907 13345 32919 13379
rect 35069 13379 35127 13385
rect 35069 13376 35081 13379
rect 32861 13339 32919 13345
rect 34164 13348 35081 13376
rect 27617 13311 27675 13317
rect 27617 13277 27629 13311
rect 27663 13277 27675 13311
rect 27617 13271 27675 13277
rect 27798 13268 27804 13320
rect 27856 13308 27862 13320
rect 29825 13311 29883 13317
rect 29825 13308 29837 13311
rect 27856 13280 29837 13308
rect 27856 13268 27862 13280
rect 29825 13277 29837 13280
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 31113 13311 31171 13317
rect 31113 13277 31125 13311
rect 31159 13277 31171 13311
rect 31113 13271 31171 13277
rect 28626 13200 28632 13252
rect 28684 13240 28690 13252
rect 28813 13243 28871 13249
rect 28813 13240 28825 13243
rect 28684 13212 28825 13240
rect 28684 13200 28690 13212
rect 28813 13209 28825 13212
rect 28859 13209 28871 13243
rect 28813 13203 28871 13209
rect 28997 13243 29055 13249
rect 28997 13209 29009 13243
rect 29043 13240 29055 13243
rect 29043 13212 30604 13240
rect 29043 13209 29055 13212
rect 28997 13203 29055 13209
rect 30466 13172 30472 13184
rect 27156 13144 30472 13172
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 30576 13172 30604 13212
rect 30742 13200 30748 13252
rect 30800 13240 30806 13252
rect 31018 13240 31024 13252
rect 30800 13212 31024 13240
rect 30800 13200 30806 13212
rect 31018 13200 31024 13212
rect 31076 13240 31082 13252
rect 31128 13240 31156 13271
rect 31202 13268 31208 13320
rect 31260 13308 31266 13320
rect 32585 13311 32643 13317
rect 32585 13308 32597 13311
rect 31260 13280 32597 13308
rect 31260 13268 31266 13280
rect 32585 13277 32597 13280
rect 32631 13277 32643 13311
rect 33870 13308 33876 13320
rect 33831 13280 33876 13308
rect 32585 13271 32643 13277
rect 33870 13268 33876 13280
rect 33928 13268 33934 13320
rect 33962 13268 33968 13320
rect 34020 13308 34026 13320
rect 34164 13317 34192 13348
rect 35069 13345 35081 13348
rect 35115 13376 35127 13379
rect 35618 13376 35624 13388
rect 35115 13348 35624 13376
rect 35115 13345 35127 13348
rect 35069 13339 35127 13345
rect 35618 13336 35624 13348
rect 35676 13336 35682 13388
rect 38102 13376 38108 13388
rect 38063 13348 38108 13376
rect 38102 13336 38108 13348
rect 38160 13336 38166 13388
rect 34149 13311 34207 13317
rect 34020 13280 34065 13308
rect 34020 13268 34026 13280
rect 34149 13277 34161 13311
rect 34195 13277 34207 13311
rect 34149 13271 34207 13277
rect 34790 13268 34796 13320
rect 34848 13308 34854 13320
rect 34885 13311 34943 13317
rect 34885 13308 34897 13311
rect 34848 13280 34897 13308
rect 34848 13268 34854 13280
rect 34885 13277 34897 13280
rect 34931 13277 34943 13311
rect 34885 13271 34943 13277
rect 35250 13268 35256 13320
rect 35308 13308 35314 13320
rect 35529 13311 35587 13317
rect 35529 13308 35541 13311
rect 35308 13280 35541 13308
rect 35308 13268 35314 13280
rect 35529 13277 35541 13280
rect 35575 13277 35587 13311
rect 35529 13271 35587 13277
rect 35986 13268 35992 13320
rect 36044 13308 36050 13320
rect 36265 13311 36323 13317
rect 36265 13308 36277 13311
rect 36044 13280 36277 13308
rect 36044 13268 36050 13280
rect 36265 13277 36277 13280
rect 36311 13277 36323 13311
rect 36265 13271 36323 13277
rect 31076 13212 31156 13240
rect 31076 13200 31082 13212
rect 35158 13200 35164 13252
rect 35216 13240 35222 13252
rect 35621 13243 35679 13249
rect 35621 13240 35633 13243
rect 35216 13212 35633 13240
rect 35216 13200 35222 13212
rect 35621 13209 35633 13212
rect 35667 13209 35679 13243
rect 35621 13203 35679 13209
rect 35805 13243 35863 13249
rect 35805 13209 35817 13243
rect 35851 13209 35863 13243
rect 35805 13203 35863 13209
rect 36449 13243 36507 13249
rect 36449 13209 36461 13243
rect 36495 13240 36507 13243
rect 37642 13240 37648 13252
rect 36495 13212 37648 13240
rect 36495 13209 36507 13212
rect 36449 13203 36507 13209
rect 31386 13172 31392 13184
rect 30576 13144 31392 13172
rect 31386 13132 31392 13144
rect 31444 13132 31450 13184
rect 34146 13132 34152 13184
rect 34204 13172 34210 13184
rect 34514 13172 34520 13184
rect 34204 13144 34520 13172
rect 34204 13132 34210 13144
rect 34514 13132 34520 13144
rect 34572 13132 34578 13184
rect 35342 13132 35348 13184
rect 35400 13172 35406 13184
rect 35706 13175 35764 13181
rect 35706 13172 35718 13175
rect 35400 13144 35718 13172
rect 35400 13132 35406 13144
rect 35706 13141 35718 13144
rect 35752 13141 35764 13175
rect 35820 13172 35848 13203
rect 37642 13200 37648 13212
rect 37700 13200 37706 13252
rect 36262 13172 36268 13184
rect 35820 13144 36268 13172
rect 35706 13135 35764 13141
rect 36262 13132 36268 13144
rect 36320 13132 36326 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 16114 12968 16120 12980
rect 15427 12940 16120 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18785 12971 18843 12977
rect 18785 12968 18797 12971
rect 18748 12940 18797 12968
rect 18748 12928 18754 12940
rect 18785 12937 18797 12940
rect 18831 12937 18843 12971
rect 19334 12968 19340 12980
rect 18785 12931 18843 12937
rect 19306 12928 19340 12968
rect 19392 12928 19398 12980
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 20772 12940 24869 12968
rect 20772 12928 20778 12940
rect 24857 12937 24869 12940
rect 24903 12968 24915 12971
rect 26418 12968 26424 12980
rect 24903 12940 26424 12968
rect 24903 12937 24915 12940
rect 24857 12931 24915 12937
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 31481 12971 31539 12977
rect 31481 12937 31493 12971
rect 31527 12968 31539 12971
rect 32283 12971 32341 12977
rect 32283 12968 32295 12971
rect 31527 12940 32295 12968
rect 31527 12937 31539 12940
rect 31481 12931 31539 12937
rect 32283 12937 32295 12940
rect 32329 12937 32341 12971
rect 32283 12931 32341 12937
rect 34054 12928 34060 12980
rect 34112 12968 34118 12980
rect 34399 12971 34457 12977
rect 34399 12968 34411 12971
rect 34112 12940 34411 12968
rect 34112 12928 34118 12940
rect 34399 12937 34411 12940
rect 34445 12937 34457 12971
rect 34399 12931 34457 12937
rect 35897 12971 35955 12977
rect 35897 12937 35909 12971
rect 35943 12968 35955 12971
rect 36446 12968 36452 12980
rect 35943 12940 36452 12968
rect 35943 12937 35955 12940
rect 35897 12931 35955 12937
rect 36446 12928 36452 12940
rect 36504 12928 36510 12980
rect 37642 12968 37648 12980
rect 37603 12940 37648 12968
rect 37642 12928 37648 12940
rect 37700 12928 37706 12980
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 14645 12903 14703 12909
rect 14645 12900 14657 12903
rect 13872 12872 14657 12900
rect 13872 12860 13878 12872
rect 14645 12869 14657 12872
rect 14691 12869 14703 12903
rect 14645 12863 14703 12869
rect 14829 12903 14887 12909
rect 14829 12869 14841 12903
rect 14875 12900 14887 12903
rect 17126 12900 17132 12912
rect 14875 12872 17132 12900
rect 14875 12869 14887 12872
rect 14829 12863 14887 12869
rect 17126 12860 17132 12872
rect 17184 12860 17190 12912
rect 19058 12900 19064 12912
rect 19019 12872 19064 12900
rect 19058 12860 19064 12872
rect 19116 12860 19122 12912
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 19208 12872 19253 12900
rect 19208 12860 19214 12872
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2958 12832 2964 12844
rect 2087 12804 2964 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2958 12792 2964 12804
rect 3016 12832 3022 12844
rect 4062 12832 4068 12844
rect 3016 12804 4068 12832
rect 3016 12792 3022 12804
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12832 14151 12835
rect 15194 12832 15200 12844
rect 14139 12804 15200 12832
rect 14139 12801 14151 12804
rect 14093 12795 14151 12801
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 16666 12832 16672 12844
rect 15611 12804 16672 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 16942 12832 16948 12844
rect 16816 12804 16948 12832
rect 16816 12792 16822 12804
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 18690 12792 18696 12844
rect 18748 12832 18754 12844
rect 19306 12841 19334 12928
rect 20990 12900 20996 12912
rect 20951 12872 20996 12900
rect 19427 12857 19485 12863
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 21174 12900 21180 12912
rect 21135 12872 21180 12900
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 22186 12900 22192 12912
rect 22112 12872 22192 12900
rect 19427 12844 19439 12857
rect 19473 12844 19485 12857
rect 18969 12835 19027 12841
rect 18969 12832 18981 12835
rect 18748 12804 18981 12832
rect 18748 12792 18754 12804
rect 18969 12801 18981 12804
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19291 12835 19349 12841
rect 19291 12801 19303 12835
rect 19337 12801 19349 12835
rect 19291 12795 19349 12801
rect 19426 12792 19432 12844
rect 19484 12792 19490 12844
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12832 20131 12835
rect 20622 12832 20628 12844
rect 20119 12804 20628 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 22112 12841 22140 12872
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 22373 12903 22431 12909
rect 22373 12869 22385 12903
rect 22419 12900 22431 12903
rect 22922 12900 22928 12912
rect 22419 12872 22928 12900
rect 22419 12869 22431 12872
rect 22373 12863 22431 12869
rect 22922 12860 22928 12872
rect 22980 12860 22986 12912
rect 23934 12900 23940 12912
rect 23308 12872 23940 12900
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12801 22155 12835
rect 22278 12832 22284 12844
rect 22239 12804 22284 12832
rect 22097 12795 22155 12801
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12832 22615 12835
rect 22646 12832 22652 12844
rect 22603 12804 22652 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 22646 12792 22652 12804
rect 22704 12792 22710 12844
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12832 22891 12835
rect 23308 12832 23336 12872
rect 23934 12860 23940 12872
rect 23992 12860 23998 12912
rect 24762 12900 24768 12912
rect 24723 12872 24768 12900
rect 24762 12860 24768 12872
rect 24820 12860 24826 12912
rect 26970 12900 26976 12912
rect 26931 12872 26976 12900
rect 26970 12860 26976 12872
rect 27028 12860 27034 12912
rect 27157 12903 27215 12909
rect 27157 12869 27169 12903
rect 27203 12900 27215 12903
rect 28626 12900 28632 12912
rect 27203 12872 28632 12900
rect 27203 12869 27215 12872
rect 27157 12863 27215 12869
rect 28626 12860 28632 12872
rect 28684 12860 28690 12912
rect 28813 12903 28871 12909
rect 28813 12869 28825 12903
rect 28859 12900 28871 12903
rect 31294 12900 31300 12912
rect 28859 12872 31300 12900
rect 28859 12869 28871 12872
rect 28813 12863 28871 12869
rect 31294 12860 31300 12872
rect 31352 12860 31358 12912
rect 32030 12900 32036 12912
rect 31404 12872 32036 12900
rect 22879 12804 23336 12832
rect 22879 12801 22891 12804
rect 22833 12795 22891 12801
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 24210 12832 24216 12844
rect 23440 12804 23485 12832
rect 24171 12804 24216 12832
rect 23440 12792 23446 12804
rect 24210 12792 24216 12804
rect 24268 12792 24274 12844
rect 25590 12832 25596 12844
rect 25551 12804 25596 12832
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 25774 12792 25780 12844
rect 25832 12832 25838 12844
rect 26237 12835 26295 12841
rect 26237 12832 26249 12835
rect 25832 12804 26249 12832
rect 25832 12792 25838 12804
rect 26237 12801 26249 12804
rect 26283 12801 26295 12835
rect 26237 12795 26295 12801
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 18782 12764 18788 12776
rect 17267 12736 18788 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 20257 12767 20315 12773
rect 20257 12733 20269 12767
rect 20303 12764 20315 12767
rect 20898 12764 20904 12776
rect 20303 12736 20904 12764
rect 20303 12733 20315 12736
rect 20257 12727 20315 12733
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 22922 12764 22928 12776
rect 21140 12736 22928 12764
rect 21140 12724 21146 12736
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 25314 12724 25320 12776
rect 25372 12764 25378 12776
rect 25409 12767 25467 12773
rect 25409 12764 25421 12767
rect 25372 12736 25421 12764
rect 25372 12724 25378 12736
rect 25409 12733 25421 12736
rect 25455 12733 25467 12767
rect 25409 12727 25467 12733
rect 25498 12724 25504 12776
rect 25556 12764 25562 12776
rect 26436 12764 26464 12795
rect 26786 12792 26792 12844
rect 26844 12832 26850 12844
rect 27893 12835 27951 12841
rect 27893 12832 27905 12835
rect 26844 12804 27905 12832
rect 26844 12792 26850 12804
rect 27893 12801 27905 12804
rect 27939 12801 27951 12835
rect 29546 12832 29552 12844
rect 29507 12804 29552 12832
rect 27893 12795 27951 12801
rect 29546 12792 29552 12804
rect 29604 12792 29610 12844
rect 29730 12832 29736 12844
rect 29691 12804 29736 12832
rect 29730 12792 29736 12804
rect 29788 12792 29794 12844
rect 29914 12832 29920 12844
rect 29875 12804 29920 12832
rect 29914 12792 29920 12804
rect 29972 12792 29978 12844
rect 30926 12792 30932 12844
rect 30984 12832 30990 12844
rect 31021 12835 31079 12841
rect 31021 12832 31033 12835
rect 30984 12804 31033 12832
rect 30984 12792 30990 12804
rect 31021 12801 31033 12804
rect 31067 12801 31079 12835
rect 31202 12832 31208 12844
rect 31163 12804 31208 12832
rect 31021 12795 31079 12801
rect 31202 12792 31208 12804
rect 31260 12792 31266 12844
rect 29638 12764 29644 12776
rect 25556 12736 26464 12764
rect 29599 12736 29644 12764
rect 25556 12724 25562 12736
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 31110 12764 31116 12776
rect 31071 12736 31116 12764
rect 31110 12724 31116 12736
rect 31168 12724 31174 12776
rect 31297 12767 31355 12773
rect 31297 12733 31309 12767
rect 31343 12764 31355 12767
rect 31404 12764 31432 12872
rect 32030 12860 32036 12872
rect 32088 12860 32094 12912
rect 32398 12860 32404 12912
rect 32456 12900 32462 12912
rect 32493 12903 32551 12909
rect 32493 12900 32505 12903
rect 32456 12872 32505 12900
rect 32456 12860 32462 12872
rect 32493 12869 32505 12872
rect 32539 12900 32551 12903
rect 33686 12900 33692 12912
rect 32539 12872 33692 12900
rect 32539 12869 32551 12872
rect 32493 12863 32551 12869
rect 33686 12860 33692 12872
rect 33744 12860 33750 12912
rect 34514 12860 34520 12912
rect 34572 12900 34578 12912
rect 34609 12903 34667 12909
rect 34609 12900 34621 12903
rect 34572 12872 34621 12900
rect 34572 12860 34578 12872
rect 34609 12869 34621 12872
rect 34655 12869 34667 12903
rect 34609 12863 34667 12869
rect 35710 12860 35716 12912
rect 35768 12900 35774 12912
rect 35768 12872 36032 12900
rect 35768 12860 35774 12872
rect 33594 12792 33600 12844
rect 33652 12832 33658 12844
rect 35342 12832 35348 12844
rect 33652 12804 35204 12832
rect 35303 12804 35348 12832
rect 33652 12792 33658 12804
rect 31343 12736 31432 12764
rect 31343 12733 31355 12736
rect 31297 12727 31355 12733
rect 19334 12656 19340 12708
rect 19392 12696 19398 12708
rect 19978 12696 19984 12708
rect 19392 12668 19984 12696
rect 19392 12656 19398 12668
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 25682 12656 25688 12708
rect 25740 12696 25746 12708
rect 30282 12696 30288 12708
rect 25740 12668 30288 12696
rect 25740 12656 25746 12668
rect 30282 12656 30288 12668
rect 30340 12656 30346 12708
rect 30374 12656 30380 12708
rect 30432 12696 30438 12708
rect 31312 12696 31340 12727
rect 32398 12724 32404 12776
rect 32456 12764 32462 12776
rect 33505 12767 33563 12773
rect 33505 12764 33517 12767
rect 32456 12736 33517 12764
rect 32456 12724 32462 12736
rect 33505 12733 33517 12736
rect 33551 12733 33563 12767
rect 33505 12727 33563 12733
rect 33781 12767 33839 12773
rect 33781 12733 33793 12767
rect 33827 12764 33839 12767
rect 33870 12764 33876 12776
rect 33827 12736 33876 12764
rect 33827 12733 33839 12736
rect 33781 12727 33839 12733
rect 33870 12724 33876 12736
rect 33928 12724 33934 12776
rect 34606 12724 34612 12776
rect 34664 12764 34670 12776
rect 35069 12767 35127 12773
rect 35069 12764 35081 12767
rect 34664 12736 35081 12764
rect 34664 12724 34670 12736
rect 35069 12733 35081 12736
rect 35115 12733 35127 12767
rect 35176 12764 35204 12804
rect 35342 12792 35348 12804
rect 35400 12792 35406 12844
rect 35802 12832 35808 12844
rect 35763 12804 35808 12832
rect 35802 12792 35808 12804
rect 35860 12792 35866 12844
rect 36004 12841 36032 12872
rect 36078 12860 36084 12912
rect 36136 12900 36142 12912
rect 36541 12903 36599 12909
rect 36541 12900 36553 12903
rect 36136 12872 36553 12900
rect 36136 12860 36142 12872
rect 36541 12869 36553 12872
rect 36587 12869 36599 12903
rect 36541 12863 36599 12869
rect 35989 12835 36047 12841
rect 35989 12801 36001 12835
rect 36035 12801 36047 12835
rect 36630 12832 36636 12844
rect 36591 12804 36636 12832
rect 35989 12795 36047 12801
rect 36630 12792 36636 12804
rect 36688 12792 36694 12844
rect 37550 12832 37556 12844
rect 37511 12804 37556 12832
rect 37550 12792 37556 12804
rect 37608 12792 37614 12844
rect 35253 12767 35311 12773
rect 35253 12764 35265 12767
rect 35176 12736 35265 12764
rect 35069 12727 35127 12733
rect 35253 12733 35265 12736
rect 35299 12733 35311 12767
rect 35253 12727 35311 12733
rect 36078 12724 36084 12776
rect 36136 12764 36142 12776
rect 36262 12764 36268 12776
rect 36136 12736 36268 12764
rect 36136 12724 36142 12736
rect 36262 12724 36268 12736
rect 36320 12724 36326 12776
rect 30432 12668 31340 12696
rect 30432 12656 30438 12668
rect 32490 12656 32496 12708
rect 32548 12696 32554 12708
rect 34241 12699 34299 12705
rect 34241 12696 34253 12699
rect 32548 12668 34253 12696
rect 32548 12656 32554 12668
rect 34241 12665 34253 12668
rect 34287 12665 34299 12699
rect 36096 12696 36124 12724
rect 34241 12659 34299 12665
rect 34440 12668 36124 12696
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1636 12600 1961 12628
rect 1636 12588 1642 12600
rect 1949 12597 1961 12600
rect 1995 12597 2007 12631
rect 13998 12628 14004 12640
rect 13959 12600 14004 12628
rect 1949 12591 2007 12597
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 23474 12628 23480 12640
rect 23435 12600 23480 12628
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 24118 12628 24124 12640
rect 24079 12600 24124 12628
rect 24118 12588 24124 12600
rect 24176 12588 24182 12640
rect 25774 12628 25780 12640
rect 25735 12600 25780 12628
rect 25774 12588 25780 12600
rect 25832 12588 25838 12640
rect 25958 12588 25964 12640
rect 26016 12628 26022 12640
rect 26329 12631 26387 12637
rect 26329 12628 26341 12631
rect 26016 12600 26341 12628
rect 26016 12588 26022 12600
rect 26329 12597 26341 12600
rect 26375 12597 26387 12631
rect 27706 12628 27712 12640
rect 27667 12600 27712 12628
rect 26329 12591 26387 12597
rect 27706 12588 27712 12600
rect 27764 12588 27770 12640
rect 29454 12628 29460 12640
rect 29415 12600 29460 12628
rect 29454 12588 29460 12600
rect 29512 12588 29518 12640
rect 31846 12588 31852 12640
rect 31904 12628 31910 12640
rect 32125 12631 32183 12637
rect 32125 12628 32137 12631
rect 31904 12600 32137 12628
rect 31904 12588 31910 12600
rect 32125 12597 32137 12600
rect 32171 12597 32183 12631
rect 32306 12628 32312 12640
rect 32267 12600 32312 12628
rect 32125 12591 32183 12597
rect 32306 12588 32312 12600
rect 32364 12588 32370 12640
rect 33962 12588 33968 12640
rect 34020 12628 34026 12640
rect 34440 12637 34468 12668
rect 34425 12631 34483 12637
rect 34425 12628 34437 12631
rect 34020 12600 34437 12628
rect 34020 12588 34026 12600
rect 34425 12597 34437 12600
rect 34471 12597 34483 12631
rect 34425 12591 34483 12597
rect 34606 12588 34612 12640
rect 34664 12628 34670 12640
rect 35161 12631 35219 12637
rect 35161 12628 35173 12631
rect 34664 12600 35173 12628
rect 34664 12588 34670 12600
rect 35161 12597 35173 12600
rect 35207 12597 35219 12631
rect 35161 12591 35219 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 18049 12427 18107 12433
rect 18049 12393 18061 12427
rect 18095 12424 18107 12427
rect 18322 12424 18328 12436
rect 18095 12396 18328 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24397 12427 24455 12433
rect 24397 12424 24409 12427
rect 24268 12396 24409 12424
rect 24268 12384 24274 12396
rect 24397 12393 24409 12396
rect 24443 12393 24455 12427
rect 24397 12387 24455 12393
rect 25590 12384 25596 12436
rect 25648 12424 25654 12436
rect 25685 12427 25743 12433
rect 25685 12424 25697 12427
rect 25648 12396 25697 12424
rect 25648 12384 25654 12396
rect 25685 12393 25697 12396
rect 25731 12393 25743 12427
rect 28810 12424 28816 12436
rect 28771 12396 28816 12424
rect 25685 12387 25743 12393
rect 28810 12384 28816 12396
rect 28868 12384 28874 12436
rect 29641 12427 29699 12433
rect 29641 12393 29653 12427
rect 29687 12424 29699 12427
rect 29730 12424 29736 12436
rect 29687 12396 29736 12424
rect 29687 12393 29699 12396
rect 29641 12387 29699 12393
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 29914 12384 29920 12436
rect 29972 12424 29978 12436
rect 31021 12427 31079 12433
rect 31021 12424 31033 12427
rect 29972 12396 31033 12424
rect 29972 12384 29978 12396
rect 31021 12393 31033 12396
rect 31067 12424 31079 12427
rect 32306 12424 32312 12436
rect 31067 12396 32312 12424
rect 31067 12393 31079 12396
rect 31021 12387 31079 12393
rect 32306 12384 32312 12396
rect 32364 12384 32370 12436
rect 33594 12384 33600 12436
rect 33652 12424 33658 12436
rect 33689 12427 33747 12433
rect 33689 12424 33701 12427
rect 33652 12396 33701 12424
rect 33652 12384 33658 12396
rect 33689 12393 33701 12396
rect 33735 12393 33747 12427
rect 33689 12387 33747 12393
rect 34422 12384 34428 12436
rect 34480 12424 34486 12436
rect 34885 12427 34943 12433
rect 34885 12424 34897 12427
rect 34480 12396 34897 12424
rect 34480 12384 34486 12396
rect 34885 12393 34897 12396
rect 34931 12393 34943 12427
rect 34885 12387 34943 12393
rect 35618 12384 35624 12436
rect 35676 12424 35682 12436
rect 35713 12427 35771 12433
rect 35713 12424 35725 12427
rect 35676 12396 35725 12424
rect 35676 12384 35682 12396
rect 35713 12393 35725 12396
rect 35759 12393 35771 12427
rect 35713 12387 35771 12393
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 21637 12359 21695 12365
rect 17092 12328 20760 12356
rect 17092 12316 17098 12328
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 1578 12288 1584 12300
rect 1539 12260 1584 12288
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 2774 12288 2780 12300
rect 2735 12260 2780 12288
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 16758 12288 16764 12300
rect 14231 12260 16764 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12288 17555 12291
rect 17954 12288 17960 12300
rect 17543 12260 17960 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 19337 12291 19395 12297
rect 19337 12288 19349 12291
rect 18748 12260 19349 12288
rect 18748 12248 18754 12260
rect 19337 12257 19349 12260
rect 19383 12257 19395 12291
rect 19337 12251 19395 12257
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12288 19855 12291
rect 20732 12288 20760 12328
rect 21637 12325 21649 12359
rect 21683 12356 21695 12359
rect 22830 12356 22836 12368
rect 21683 12328 22836 12356
rect 21683 12325 21695 12328
rect 21637 12319 21695 12325
rect 22830 12316 22836 12328
rect 22888 12316 22894 12368
rect 30469 12359 30527 12365
rect 30469 12325 30481 12359
rect 30515 12356 30527 12359
rect 30515 12328 32260 12356
rect 30515 12325 30527 12328
rect 30469 12319 30527 12325
rect 23474 12288 23480 12300
rect 19843 12260 20668 12288
rect 20732 12260 23480 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 17221 12223 17279 12229
rect 15988 12192 16033 12220
rect 15988 12180 15994 12192
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 18046 12220 18052 12232
rect 17267 12192 18052 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 18046 12180 18052 12192
rect 18104 12220 18110 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 18104 12192 18245 12220
rect 18104 12180 18110 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12220 18475 12223
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 18463 12192 19441 12220
rect 18463 12189 18475 12192
rect 18417 12183 18475 12189
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 15657 12155 15715 12161
rect 14056 12124 14490 12152
rect 14056 12112 14062 12124
rect 15657 12121 15669 12155
rect 15703 12152 15715 12155
rect 18601 12155 18659 12161
rect 15703 12124 18552 12152
rect 15703 12121 15715 12124
rect 15657 12115 15715 12121
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 16853 12087 16911 12093
rect 16853 12084 16865 12087
rect 14424 12056 16865 12084
rect 14424 12044 14430 12056
rect 16853 12053 16865 12056
rect 16899 12053 16911 12087
rect 16853 12047 16911 12053
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17368 12056 17413 12084
rect 17368 12044 17374 12056
rect 17770 12044 17776 12096
rect 17828 12084 17834 12096
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 17828 12056 18337 12084
rect 17828 12044 17834 12056
rect 18325 12053 18337 12056
rect 18371 12053 18383 12087
rect 18524 12084 18552 12124
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 18782 12152 18788 12164
rect 18647 12124 18788 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 19242 12112 19248 12164
rect 19300 12152 19306 12164
rect 19444 12152 19472 12183
rect 20070 12180 20076 12232
rect 20128 12220 20134 12232
rect 20640 12229 20668 12260
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 25041 12291 25099 12297
rect 25041 12257 25053 12291
rect 25087 12288 25099 12291
rect 25958 12288 25964 12300
rect 25087 12260 25964 12288
rect 25087 12257 25099 12260
rect 25041 12251 25099 12257
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 32232 12297 32260 12328
rect 32217 12291 32275 12297
rect 32217 12257 32229 12291
rect 32263 12257 32275 12291
rect 32398 12288 32404 12300
rect 32359 12260 32404 12288
rect 32217 12251 32275 12257
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 20128 12192 20453 12220
rect 20128 12180 20134 12192
rect 20441 12189 20453 12192
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12220 20867 12223
rect 20898 12220 20904 12232
rect 20855 12192 20904 12220
rect 20855 12189 20867 12192
rect 20809 12183 20867 12189
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 21545 12223 21603 12229
rect 21545 12220 21557 12223
rect 21232 12192 21557 12220
rect 21232 12180 21238 12192
rect 21545 12189 21557 12192
rect 21591 12189 21603 12223
rect 21910 12220 21916 12232
rect 21871 12192 21916 12220
rect 21545 12183 21603 12189
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 22370 12220 22376 12232
rect 22331 12192 22376 12220
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22922 12180 22928 12232
rect 22980 12220 22986 12232
rect 23017 12223 23075 12229
rect 23017 12220 23029 12223
rect 22980 12192 23029 12220
rect 22980 12180 22986 12192
rect 23017 12189 23029 12192
rect 23063 12189 23075 12223
rect 23492 12220 23520 12248
rect 23661 12223 23719 12229
rect 23661 12220 23673 12223
rect 23492 12192 23673 12220
rect 23017 12183 23075 12189
rect 23661 12189 23673 12192
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12220 23903 12223
rect 24762 12220 24768 12232
rect 23891 12192 24768 12220
rect 23891 12189 23903 12192
rect 23845 12183 23903 12189
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 25406 12180 25412 12232
rect 25464 12220 25470 12232
rect 25593 12223 25651 12229
rect 25593 12220 25605 12223
rect 25464 12192 25605 12220
rect 25464 12180 25470 12192
rect 25593 12189 25605 12192
rect 25639 12189 25651 12223
rect 25593 12183 25651 12189
rect 25869 12223 25927 12229
rect 25869 12189 25881 12223
rect 25915 12220 25927 12223
rect 26326 12220 26332 12232
rect 25915 12192 26332 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 26326 12180 26332 12192
rect 26384 12180 26390 12232
rect 26602 12220 26608 12232
rect 26563 12192 26608 12220
rect 26602 12180 26608 12192
rect 26660 12180 26666 12232
rect 28994 12220 29000 12232
rect 28955 12192 29000 12220
rect 28994 12180 29000 12192
rect 29052 12180 29058 12232
rect 29733 12223 29791 12229
rect 29733 12189 29745 12223
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 30193 12223 30251 12229
rect 30193 12189 30205 12223
rect 30239 12220 30251 12223
rect 30374 12220 30380 12232
rect 30239 12192 30380 12220
rect 30239 12189 30251 12192
rect 30193 12183 30251 12189
rect 20533 12155 20591 12161
rect 20533 12152 20545 12155
rect 19300 12124 20545 12152
rect 19300 12112 19306 12124
rect 20533 12121 20545 12124
rect 20579 12121 20591 12155
rect 23201 12155 23259 12161
rect 23201 12152 23213 12155
rect 20533 12115 20591 12121
rect 22066 12124 23213 12152
rect 20257 12087 20315 12093
rect 20257 12084 20269 12087
rect 18524 12056 20269 12084
rect 18325 12047 18383 12053
rect 20257 12053 20269 12056
rect 20303 12053 20315 12087
rect 20257 12047 20315 12053
rect 20622 12044 20628 12096
rect 20680 12084 20686 12096
rect 22066 12084 22094 12124
rect 23201 12121 23213 12124
rect 23247 12152 23259 12155
rect 23566 12152 23572 12164
rect 23247 12124 23572 12152
rect 23247 12121 23259 12124
rect 23201 12115 23259 12121
rect 23566 12112 23572 12124
rect 23624 12112 23630 12164
rect 23753 12155 23811 12161
rect 23753 12121 23765 12155
rect 23799 12152 23811 12155
rect 24857 12155 24915 12161
rect 24857 12152 24869 12155
rect 23799 12124 24869 12152
rect 23799 12121 23811 12124
rect 23753 12115 23811 12121
rect 24857 12121 24869 12124
rect 24903 12121 24915 12155
rect 24857 12115 24915 12121
rect 26053 12155 26111 12161
rect 26053 12121 26065 12155
rect 26099 12152 26111 12155
rect 26881 12155 26939 12161
rect 26881 12152 26893 12155
rect 26099 12124 26893 12152
rect 26099 12121 26111 12124
rect 26053 12115 26111 12121
rect 26881 12121 26893 12124
rect 26927 12121 26939 12155
rect 26881 12115 26939 12121
rect 27614 12112 27620 12164
rect 27672 12112 27678 12164
rect 29748 12152 29776 12183
rect 30374 12180 30380 12192
rect 30432 12180 30438 12232
rect 30466 12180 30472 12232
rect 30524 12220 30530 12232
rect 30926 12220 30932 12232
rect 30524 12192 30569 12220
rect 30887 12192 30932 12220
rect 30524 12180 30530 12192
rect 30926 12180 30932 12192
rect 30984 12180 30990 12232
rect 31018 12180 31024 12232
rect 31076 12220 31082 12232
rect 31297 12223 31355 12229
rect 31297 12220 31309 12223
rect 31076 12192 31309 12220
rect 31076 12180 31082 12192
rect 31297 12189 31309 12192
rect 31343 12189 31355 12223
rect 32232 12220 32260 12251
rect 32398 12248 32404 12260
rect 32456 12248 32462 12300
rect 36814 12288 36820 12300
rect 35820 12260 36820 12288
rect 33505 12223 33563 12229
rect 33505 12220 33517 12223
rect 32232 12192 33517 12220
rect 31297 12183 31355 12189
rect 33505 12189 33517 12192
rect 33551 12189 33563 12223
rect 33505 12183 33563 12189
rect 33781 12223 33839 12229
rect 33781 12189 33793 12223
rect 33827 12220 33839 12223
rect 34146 12220 34152 12232
rect 33827 12192 34152 12220
rect 33827 12189 33839 12192
rect 33781 12183 33839 12189
rect 34146 12180 34152 12192
rect 34204 12180 34210 12232
rect 35820 12229 35848 12260
rect 36814 12248 36820 12260
rect 36872 12248 36878 12300
rect 34977 12223 35035 12229
rect 34977 12189 34989 12223
rect 35023 12220 35035 12223
rect 35805 12223 35863 12229
rect 35805 12220 35817 12223
rect 35023 12192 35817 12220
rect 35023 12189 35035 12192
rect 34977 12183 35035 12189
rect 35805 12189 35817 12192
rect 35851 12189 35863 12223
rect 36262 12220 36268 12232
rect 36223 12192 36268 12220
rect 35805 12183 35863 12189
rect 36262 12180 36268 12192
rect 36320 12180 36326 12232
rect 30742 12152 30748 12164
rect 29748 12124 30748 12152
rect 30742 12112 30748 12124
rect 30800 12112 30806 12164
rect 31202 12152 31208 12164
rect 30944 12124 31208 12152
rect 24762 12084 24768 12096
rect 20680 12056 22094 12084
rect 24723 12056 24768 12084
rect 20680 12044 20686 12056
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 28353 12087 28411 12093
rect 28353 12053 28365 12087
rect 28399 12084 28411 12087
rect 29362 12084 29368 12096
rect 28399 12056 29368 12084
rect 28399 12053 28411 12056
rect 28353 12047 28411 12053
rect 29362 12044 29368 12056
rect 29420 12044 29426 12096
rect 30285 12087 30343 12093
rect 30285 12053 30297 12087
rect 30331 12084 30343 12087
rect 30944 12084 30972 12124
rect 31202 12112 31208 12124
rect 31260 12112 31266 12164
rect 32398 12152 32404 12164
rect 31312 12124 32404 12152
rect 31110 12084 31116 12096
rect 30331 12056 30972 12084
rect 31023 12056 31116 12084
rect 30331 12053 30343 12056
rect 30285 12047 30343 12053
rect 31110 12044 31116 12056
rect 31168 12084 31174 12096
rect 31312 12084 31340 12124
rect 32398 12112 32404 12124
rect 32456 12112 32462 12164
rect 36449 12155 36507 12161
rect 36449 12121 36461 12155
rect 36495 12152 36507 12155
rect 37642 12152 37648 12164
rect 36495 12124 37648 12152
rect 36495 12121 36507 12124
rect 36449 12115 36507 12121
rect 37642 12112 37648 12124
rect 37700 12112 37706 12164
rect 38102 12152 38108 12164
rect 38063 12124 38108 12152
rect 38102 12112 38108 12124
rect 38160 12112 38166 12164
rect 31754 12084 31760 12096
rect 31168 12056 31340 12084
rect 31715 12056 31760 12084
rect 31168 12044 31174 12056
rect 31754 12044 31760 12056
rect 31812 12044 31818 12096
rect 32122 12084 32128 12096
rect 32083 12056 32128 12084
rect 32122 12044 32128 12056
rect 32180 12044 32186 12096
rect 32674 12044 32680 12096
rect 32732 12084 32738 12096
rect 33321 12087 33379 12093
rect 33321 12084 33333 12087
rect 32732 12056 33333 12084
rect 32732 12044 32738 12056
rect 33321 12053 33333 12056
rect 33367 12053 33379 12087
rect 33321 12047 33379 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 13078 11880 13084 11892
rect 12912 11852 13084 11880
rect 12912 11753 12940 11852
rect 13078 11840 13084 11852
rect 13136 11880 13142 11892
rect 13906 11880 13912 11892
rect 13136 11852 13912 11880
rect 13136 11840 13142 11852
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 17221 11883 17279 11889
rect 17221 11849 17233 11883
rect 17267 11880 17279 11883
rect 17310 11880 17316 11892
rect 17267 11852 17316 11880
rect 17267 11849 17279 11852
rect 17221 11843 17279 11849
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 17552 11852 17693 11880
rect 17552 11840 17558 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 17681 11843 17739 11849
rect 17849 11883 17907 11889
rect 17849 11849 17861 11883
rect 17895 11880 17907 11883
rect 17954 11880 17960 11892
rect 17895 11852 17960 11880
rect 17895 11849 17907 11852
rect 17849 11843 17907 11849
rect 17954 11840 17960 11852
rect 18012 11880 18018 11892
rect 18230 11880 18236 11892
rect 18012 11852 18236 11880
rect 18012 11840 18018 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 18598 11880 18604 11892
rect 18559 11852 18604 11880
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 20622 11880 20628 11892
rect 19076 11852 20628 11880
rect 19076 11824 19104 11852
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 21269 11883 21327 11889
rect 21269 11849 21281 11883
rect 21315 11880 21327 11883
rect 21910 11880 21916 11892
rect 21315 11852 21916 11880
rect 21315 11849 21327 11852
rect 21269 11843 21327 11849
rect 21910 11840 21916 11852
rect 21968 11840 21974 11892
rect 25774 11880 25780 11892
rect 25735 11852 25780 11880
rect 25774 11840 25780 11852
rect 25832 11840 25838 11892
rect 26145 11883 26203 11889
rect 26145 11849 26157 11883
rect 26191 11880 26203 11883
rect 26786 11880 26792 11892
rect 26191 11852 26792 11880
rect 26191 11849 26203 11852
rect 26145 11843 26203 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 30466 11880 30472 11892
rect 29288 11852 30472 11880
rect 15194 11772 15200 11824
rect 15252 11812 15258 11824
rect 15381 11815 15439 11821
rect 15381 11812 15393 11815
rect 15252 11784 15393 11812
rect 15252 11772 15258 11784
rect 15381 11781 15393 11784
rect 15427 11781 15439 11815
rect 15381 11775 15439 11781
rect 18049 11815 18107 11821
rect 18049 11781 18061 11815
rect 18095 11812 18107 11815
rect 19058 11812 19064 11824
rect 18095 11784 19064 11812
rect 18095 11781 18107 11784
rect 18049 11775 18107 11781
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 20438 11772 20444 11824
rect 20496 11812 20502 11824
rect 22005 11815 22063 11821
rect 22005 11812 22017 11815
rect 20496 11784 22017 11812
rect 20496 11772 20502 11784
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 14274 11704 14280 11756
rect 14332 11704 14338 11756
rect 15562 11744 15568 11756
rect 15475 11716 15568 11744
rect 15562 11704 15568 11716
rect 15620 11744 15626 11756
rect 16114 11744 16120 11756
rect 15620 11716 16120 11744
rect 15620 11704 15626 11716
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 18509 11747 18567 11753
rect 17267 11716 18092 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 18064 11688 18092 11716
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 18690 11744 18696 11756
rect 18651 11716 18696 11744
rect 18509 11707 18567 11713
rect 1578 11676 1584 11688
rect 1539 11648 1584 11676
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 1946 11676 1952 11688
rect 1811 11648 1952 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 13173 11679 13231 11685
rect 2096 11648 2141 11676
rect 2096 11636 2102 11648
rect 13173 11645 13185 11679
rect 13219 11676 13231 11679
rect 14182 11676 14188 11688
rect 13219 11648 14188 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 18524 11676 18552 11707
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19300 11716 19809 11744
rect 19300 11704 19306 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 19978 11704 19984 11756
rect 20036 11744 20042 11756
rect 21100 11753 21128 11784
rect 22005 11781 22017 11784
rect 22051 11781 22063 11815
rect 24670 11812 24676 11824
rect 24334 11784 24676 11812
rect 22005 11775 22063 11781
rect 24670 11772 24676 11784
rect 24728 11772 24734 11824
rect 25685 11815 25743 11821
rect 25685 11781 25697 11815
rect 25731 11812 25743 11815
rect 26326 11812 26332 11824
rect 25731 11784 26332 11812
rect 25731 11781 25743 11784
rect 25685 11775 25743 11781
rect 26326 11772 26332 11784
rect 26384 11772 26390 11824
rect 29288 11812 29316 11852
rect 30466 11840 30472 11852
rect 30524 11840 30530 11892
rect 30742 11840 30748 11892
rect 30800 11880 30806 11892
rect 30929 11883 30987 11889
rect 30929 11880 30941 11883
rect 30800 11852 30941 11880
rect 30800 11840 30806 11852
rect 30929 11849 30941 11852
rect 30975 11880 30987 11883
rect 31570 11880 31576 11892
rect 30975 11852 31576 11880
rect 30975 11849 30987 11852
rect 30929 11843 30987 11849
rect 31570 11840 31576 11852
rect 31628 11840 31634 11892
rect 32122 11880 32128 11892
rect 32083 11852 32128 11880
rect 32122 11840 32128 11852
rect 32180 11840 32186 11892
rect 36078 11880 36084 11892
rect 36039 11852 36084 11880
rect 36078 11840 36084 11852
rect 36136 11840 36142 11892
rect 37642 11880 37648 11892
rect 37603 11852 37648 11880
rect 37642 11840 37648 11852
rect 37700 11840 37706 11892
rect 29454 11812 29460 11824
rect 28474 11784 29316 11812
rect 29415 11784 29460 11812
rect 29454 11772 29460 11784
rect 29512 11772 29518 11824
rect 29914 11772 29920 11824
rect 29972 11772 29978 11824
rect 32030 11772 32036 11824
rect 32088 11812 32094 11824
rect 32277 11815 32335 11821
rect 32277 11812 32289 11815
rect 32088 11784 32289 11812
rect 32088 11772 32094 11784
rect 32277 11781 32289 11784
rect 32323 11781 32335 11815
rect 32490 11812 32496 11824
rect 32451 11784 32496 11812
rect 32277 11775 32335 11781
rect 32490 11772 32496 11784
rect 32548 11772 32554 11824
rect 34606 11812 34612 11824
rect 34567 11784 34612 11812
rect 34606 11772 34612 11784
rect 34664 11772 34670 11824
rect 35342 11772 35348 11824
rect 35400 11772 35406 11824
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 20036 11716 20821 11744
rect 20036 11704 20042 11716
rect 20809 11713 20821 11716
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 21821 11747 21879 11753
rect 21821 11713 21833 11747
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 31389 11747 31447 11753
rect 31389 11713 31401 11747
rect 31435 11744 31447 11747
rect 31846 11744 31852 11756
rect 31435 11716 31852 11744
rect 31435 11713 31447 11716
rect 31389 11707 31447 11713
rect 19260 11676 19288 11704
rect 18524 11648 19288 11676
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 19484 11648 20085 11676
rect 19484 11636 19490 11648
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 20993 11679 21051 11685
rect 20993 11645 21005 11679
rect 21039 11676 21051 11679
rect 21450 11676 21456 11688
rect 21039 11648 21456 11676
rect 21039 11645 21051 11648
rect 20993 11639 21051 11645
rect 21450 11636 21456 11648
rect 21508 11636 21514 11688
rect 21836 11608 21864 11707
rect 31846 11704 31852 11716
rect 31904 11704 31910 11756
rect 32950 11744 32956 11756
rect 32911 11716 32956 11744
rect 32950 11704 32956 11716
rect 33008 11704 33014 11756
rect 36722 11744 36728 11756
rect 36635 11716 36728 11744
rect 36722 11704 36728 11716
rect 36780 11744 36786 11756
rect 37734 11744 37740 11756
rect 36780 11716 37740 11744
rect 36780 11704 36786 11716
rect 37734 11704 37740 11716
rect 37792 11704 37798 11756
rect 22833 11679 22891 11685
rect 22833 11645 22845 11679
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 23109 11679 23167 11685
rect 23109 11645 23121 11679
rect 23155 11676 23167 11679
rect 24118 11676 24124 11688
rect 23155 11648 24124 11676
rect 23155 11645 23167 11648
rect 23109 11639 23167 11645
rect 20824 11580 21864 11608
rect 14645 11543 14703 11549
rect 14645 11509 14657 11543
rect 14691 11540 14703 11543
rect 16850 11540 16856 11552
rect 14691 11512 16856 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17865 11543 17923 11549
rect 17865 11509 17877 11543
rect 17911 11540 17923 11543
rect 18322 11540 18328 11552
rect 17911 11512 18328 11540
rect 17911 11509 17923 11512
rect 17865 11503 17923 11509
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 18598 11500 18604 11552
rect 18656 11540 18662 11552
rect 20070 11540 20076 11552
rect 18656 11512 20076 11540
rect 18656 11500 18662 11512
rect 20070 11500 20076 11512
rect 20128 11540 20134 11552
rect 20438 11540 20444 11552
rect 20128 11512 20444 11540
rect 20128 11500 20134 11512
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 20824 11549 20852 11580
rect 20809 11543 20867 11549
rect 20809 11540 20821 11543
rect 20588 11512 20821 11540
rect 20588 11500 20594 11512
rect 20809 11509 20821 11512
rect 20855 11509 20867 11543
rect 20809 11503 20867 11509
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22189 11543 22247 11549
rect 22189 11540 22201 11543
rect 22152 11512 22201 11540
rect 22152 11500 22158 11512
rect 22189 11509 22201 11512
rect 22235 11509 22247 11543
rect 22189 11503 22247 11509
rect 22462 11500 22468 11552
rect 22520 11540 22526 11552
rect 22646 11540 22652 11552
rect 22520 11512 22652 11540
rect 22520 11500 22526 11512
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 22848 11540 22876 11639
rect 24118 11636 24124 11648
rect 24176 11636 24182 11688
rect 25590 11676 25596 11688
rect 25551 11648 25596 11676
rect 25590 11636 25596 11648
rect 25648 11636 25654 11688
rect 26973 11679 27031 11685
rect 26973 11645 26985 11679
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 27249 11679 27307 11685
rect 27249 11645 27261 11679
rect 27295 11676 27307 11679
rect 27706 11676 27712 11688
rect 27295 11648 27712 11676
rect 27295 11645 27307 11648
rect 27249 11639 27307 11645
rect 26234 11608 26240 11620
rect 24136 11580 26240 11608
rect 24136 11540 24164 11580
rect 26234 11568 26240 11580
rect 26292 11608 26298 11620
rect 26602 11608 26608 11620
rect 26292 11580 26608 11608
rect 26292 11568 26298 11580
rect 26602 11568 26608 11580
rect 26660 11608 26666 11620
rect 26988 11608 27016 11639
rect 27706 11636 27712 11648
rect 27764 11636 27770 11688
rect 28718 11636 28724 11688
rect 28776 11676 28782 11688
rect 29181 11679 29239 11685
rect 29181 11676 29193 11679
rect 28776 11648 29193 11676
rect 28776 11636 28782 11648
rect 29181 11645 29193 11648
rect 29227 11645 29239 11679
rect 29181 11639 29239 11645
rect 26660 11580 27016 11608
rect 26660 11568 26666 11580
rect 24578 11540 24584 11552
rect 22848 11512 24164 11540
rect 24539 11512 24584 11540
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 28626 11500 28632 11552
rect 28684 11540 28690 11552
rect 28721 11543 28779 11549
rect 28721 11540 28733 11543
rect 28684 11512 28733 11540
rect 28684 11500 28690 11512
rect 28721 11509 28733 11512
rect 28767 11509 28779 11543
rect 29196 11540 29224 11639
rect 31662 11636 31668 11688
rect 31720 11676 31726 11688
rect 34333 11679 34391 11685
rect 34333 11676 34345 11679
rect 31720 11648 34345 11676
rect 31720 11636 31726 11648
rect 34333 11645 34345 11648
rect 34379 11645 34391 11679
rect 34333 11639 34391 11645
rect 31202 11568 31208 11620
rect 31260 11608 31266 11620
rect 31260 11580 32352 11608
rect 31260 11568 31266 11580
rect 30834 11540 30840 11552
rect 29196 11512 30840 11540
rect 28721 11503 28779 11509
rect 30834 11500 30840 11512
rect 30892 11500 30898 11552
rect 31570 11540 31576 11552
rect 31531 11512 31576 11540
rect 31570 11500 31576 11512
rect 31628 11500 31634 11552
rect 32324 11549 32352 11580
rect 32309 11543 32367 11549
rect 32309 11509 32321 11543
rect 32355 11509 32367 11543
rect 32309 11503 32367 11509
rect 33045 11543 33103 11549
rect 33045 11509 33057 11543
rect 33091 11540 33103 11543
rect 33410 11540 33416 11552
rect 33091 11512 33416 11540
rect 33091 11509 33103 11512
rect 33045 11503 33103 11509
rect 33410 11500 33416 11512
rect 33468 11500 33474 11552
rect 33873 11543 33931 11549
rect 33873 11509 33885 11543
rect 33919 11540 33931 11543
rect 35894 11540 35900 11552
rect 33919 11512 35900 11540
rect 33919 11509 33931 11512
rect 33873 11503 33931 11509
rect 35894 11500 35900 11512
rect 35952 11500 35958 11552
rect 36538 11500 36544 11552
rect 36596 11540 36602 11552
rect 36633 11543 36691 11549
rect 36633 11540 36645 11543
rect 36596 11512 36645 11540
rect 36596 11500 36602 11512
rect 36633 11509 36645 11512
rect 36679 11509 36691 11543
rect 36633 11503 36691 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 14182 11336 14188 11348
rect 14143 11308 14188 11336
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 17310 11336 17316 11348
rect 14967 11308 17316 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 17589 11339 17647 11345
rect 17589 11305 17601 11339
rect 17635 11336 17647 11339
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 17635 11308 19441 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 22462 11296 22468 11348
rect 22520 11336 22526 11348
rect 22649 11339 22707 11345
rect 22649 11336 22661 11339
rect 22520 11308 22661 11336
rect 22520 11296 22526 11308
rect 22649 11305 22661 11308
rect 22695 11305 22707 11339
rect 22649 11299 22707 11305
rect 22922 11296 22928 11348
rect 22980 11336 22986 11348
rect 22980 11308 26188 11336
rect 22980 11296 22986 11308
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 18708 11240 19257 11268
rect 15930 11160 15936 11212
rect 15988 11200 15994 11212
rect 16390 11200 16396 11212
rect 15988 11172 16396 11200
rect 15988 11160 15994 11172
rect 16390 11160 16396 11172
rect 16448 11200 16454 11212
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 16448 11172 16681 11200
rect 16448 11160 16454 11172
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 17954 11200 17960 11212
rect 16669 11163 16727 11169
rect 17328 11172 17960 11200
rect 2038 11132 2044 11144
rect 1951 11104 2044 11132
rect 2038 11092 2044 11104
rect 2096 11132 2102 11144
rect 2222 11132 2228 11144
rect 2096 11104 2228 11132
rect 2096 11092 2102 11104
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14366 11132 14372 11144
rect 14323 11104 14372 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 17328 11141 17356 11172
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11200 18291 11203
rect 18598 11200 18604 11212
rect 18279 11172 18604 11200
rect 18279 11169 18291 11172
rect 18233 11163 18291 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 18708 11209 18736 11240
rect 19245 11237 19257 11240
rect 19291 11237 19303 11271
rect 19245 11231 19303 11237
rect 21100 11240 22094 11268
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11169 18751 11203
rect 18693 11163 18751 11169
rect 19168 11172 20760 11200
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11101 17371 11135
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 17313 11095 17371 11101
rect 17420 11104 18061 11132
rect 16393 11067 16451 11073
rect 16393 11033 16405 11067
rect 16439 11064 16451 11067
rect 17420 11064 17448 11104
rect 18049 11101 18061 11104
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 19168 11132 19196 11172
rect 18371 11104 19196 11132
rect 19429 11135 19487 11141
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 20254 11132 20260 11144
rect 19659 11104 20260 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 16439 11036 17448 11064
rect 17589 11067 17647 11073
rect 16439 11033 16451 11036
rect 16393 11027 16451 11033
rect 17589 11033 17601 11067
rect 17635 11064 17647 11067
rect 17770 11064 17776 11076
rect 17635 11036 17776 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 17770 11024 17776 11036
rect 17828 11064 17834 11076
rect 18340 11064 18368 11095
rect 17828 11036 18368 11064
rect 17828 11024 17834 11036
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 19444 11064 19472 11095
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 20732 11141 20760 11172
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11132 20775 11135
rect 20898 11132 20904 11144
rect 20763 11104 20904 11132
rect 20763 11101 20775 11104
rect 20717 11095 20775 11101
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11132 21051 11135
rect 21100 11132 21128 11240
rect 21450 11200 21456 11212
rect 21411 11172 21456 11200
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 21039 11104 21128 11132
rect 21039 11101 21051 11104
rect 20993 11095 21051 11101
rect 18748 11036 19472 11064
rect 18748 11024 18754 11036
rect 20070 11024 20076 11076
rect 20128 11064 20134 11076
rect 21008 11064 21036 11095
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 21652 11141 21864 11142
rect 21652 11135 21879 11141
rect 21652 11132 21833 11135
rect 21600 11114 21833 11132
rect 21600 11104 21680 11114
rect 21600 11092 21606 11104
rect 21821 11101 21833 11114
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 21949 11135 22007 11141
rect 21949 11101 21961 11135
rect 21995 11132 22007 11135
rect 22066 11132 22094 11240
rect 24118 11228 24124 11280
rect 24176 11268 24182 11280
rect 24762 11268 24768 11280
rect 24176 11240 24768 11268
rect 24176 11228 24182 11240
rect 22833 11203 22891 11209
rect 22833 11169 22845 11203
rect 22879 11200 22891 11203
rect 23750 11200 23756 11212
rect 22879 11172 23756 11200
rect 22879 11169 22891 11172
rect 22833 11163 22891 11169
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 24397 11203 24455 11209
rect 24397 11169 24409 11203
rect 24443 11200 24455 11203
rect 24578 11200 24584 11212
rect 24443 11172 24584 11200
rect 24443 11169 24455 11172
rect 24397 11163 24455 11169
rect 24578 11160 24584 11172
rect 24636 11160 24642 11212
rect 24688 11209 24716 11240
rect 24762 11228 24768 11240
rect 24820 11228 24826 11280
rect 25222 11228 25228 11280
rect 25280 11268 25286 11280
rect 26160 11268 26188 11308
rect 26694 11296 26700 11348
rect 26752 11336 26758 11348
rect 26789 11339 26847 11345
rect 26789 11336 26801 11339
rect 26752 11308 26801 11336
rect 26752 11296 26758 11308
rect 26789 11305 26801 11308
rect 26835 11305 26847 11339
rect 26789 11299 26847 11305
rect 27430 11296 27436 11348
rect 27488 11336 27494 11348
rect 27525 11339 27583 11345
rect 27525 11336 27537 11339
rect 27488 11308 27537 11336
rect 27488 11296 27494 11308
rect 27525 11305 27537 11308
rect 27571 11305 27583 11339
rect 27525 11299 27583 11305
rect 29641 11339 29699 11345
rect 29641 11305 29653 11339
rect 29687 11336 29699 11339
rect 29914 11336 29920 11348
rect 29687 11308 29920 11336
rect 29687 11305 29699 11308
rect 29641 11299 29699 11305
rect 29914 11296 29920 11308
rect 29972 11296 29978 11348
rect 30193 11339 30251 11345
rect 30193 11305 30205 11339
rect 30239 11336 30251 11339
rect 30926 11336 30932 11348
rect 30239 11308 30932 11336
rect 30239 11305 30251 11308
rect 30193 11299 30251 11305
rect 30926 11296 30932 11308
rect 30984 11296 30990 11348
rect 34146 11336 34152 11348
rect 34107 11308 34152 11336
rect 34146 11296 34152 11308
rect 34204 11296 34210 11348
rect 35069 11339 35127 11345
rect 35069 11305 35081 11339
rect 35115 11336 35127 11339
rect 35434 11336 35440 11348
rect 35115 11308 35440 11336
rect 35115 11305 35127 11308
rect 35069 11299 35127 11305
rect 35434 11296 35440 11308
rect 35492 11296 35498 11348
rect 29178 11268 29184 11280
rect 25280 11240 26096 11268
rect 26160 11240 29184 11268
rect 25280 11228 25286 11240
rect 26068 11212 26096 11240
rect 29178 11228 29184 11240
rect 29236 11228 29242 11280
rect 34698 11228 34704 11280
rect 34756 11268 34762 11280
rect 35713 11271 35771 11277
rect 35713 11268 35725 11271
rect 34756 11240 35725 11268
rect 34756 11228 34762 11240
rect 35713 11237 35725 11240
rect 35759 11237 35771 11271
rect 35713 11231 35771 11237
rect 36078 11228 36084 11280
rect 36136 11268 36142 11280
rect 36814 11268 36820 11280
rect 36136 11240 36820 11268
rect 36136 11228 36142 11240
rect 36814 11228 36820 11240
rect 36872 11228 36878 11280
rect 24673 11203 24731 11209
rect 24673 11169 24685 11203
rect 24719 11169 24731 11203
rect 24673 11163 24731 11169
rect 25314 11160 25320 11212
rect 25372 11200 25378 11212
rect 25685 11203 25743 11209
rect 25685 11200 25697 11203
rect 25372 11172 25697 11200
rect 25372 11160 25378 11172
rect 25685 11169 25697 11172
rect 25731 11169 25743 11203
rect 26050 11200 26056 11212
rect 25963 11172 26056 11200
rect 25685 11163 25743 11169
rect 26050 11160 26056 11172
rect 26108 11160 26114 11212
rect 27246 11200 27252 11212
rect 26896 11172 27252 11200
rect 21995 11104 22094 11132
rect 22649 11135 22707 11141
rect 21995 11101 22007 11104
rect 21949 11095 22007 11101
rect 22649 11101 22661 11135
rect 22695 11132 22707 11135
rect 22695 11104 22876 11132
rect 22695 11101 22707 11104
rect 22649 11095 22707 11101
rect 21637 11067 21695 11073
rect 21637 11064 21649 11067
rect 20128 11036 21036 11064
rect 21100 11036 21649 11064
rect 20128 11024 20134 11036
rect 17405 10999 17463 11005
rect 17405 10965 17417 10999
rect 17451 10996 17463 10999
rect 18046 10996 18052 11008
rect 17451 10968 18052 10996
rect 17451 10965 17463 10968
rect 17405 10959 17463 10965
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 20806 10956 20812 11008
rect 20864 10996 20870 11008
rect 21100 10996 21128 11036
rect 21637 11033 21649 11036
rect 21683 11033 21695 11067
rect 21637 11027 21695 11033
rect 21729 11067 21787 11073
rect 21729 11033 21741 11067
rect 21775 11033 21787 11067
rect 22848 11064 22876 11104
rect 22922 11092 22928 11144
rect 22980 11132 22986 11144
rect 23566 11132 23572 11144
rect 22980 11104 23025 11132
rect 23479 11104 23572 11132
rect 22980 11092 22986 11104
rect 23566 11092 23572 11104
rect 23624 11132 23630 11144
rect 24026 11132 24032 11144
rect 23624 11104 24032 11132
rect 23624 11092 23630 11104
rect 24026 11092 24032 11104
rect 24084 11092 24090 11144
rect 24302 11092 24308 11144
rect 24360 11132 24366 11144
rect 25869 11135 25927 11141
rect 25869 11132 25881 11135
rect 24360 11104 25881 11132
rect 24360 11092 24366 11104
rect 25869 11101 25881 11104
rect 25915 11101 25927 11135
rect 25869 11095 25927 11101
rect 25958 11092 25964 11144
rect 26016 11132 26022 11144
rect 26145 11135 26203 11141
rect 26016 11104 26061 11132
rect 26016 11092 26022 11104
rect 26145 11101 26157 11135
rect 26191 11132 26203 11135
rect 26694 11132 26700 11144
rect 26191 11104 26700 11132
rect 26191 11101 26203 11104
rect 26145 11095 26203 11101
rect 23842 11064 23848 11076
rect 21729 11027 21787 11033
rect 22112 11036 22784 11064
rect 22848 11036 23848 11064
rect 20864 10968 21128 10996
rect 21744 10996 21772 11027
rect 22112 10996 22140 11036
rect 21744 10968 22140 10996
rect 20864 10956 20870 10968
rect 22186 10956 22192 11008
rect 22244 10996 22250 11008
rect 22465 10999 22523 11005
rect 22465 10996 22477 10999
rect 22244 10968 22477 10996
rect 22244 10956 22250 10968
rect 22465 10965 22477 10968
rect 22511 10965 22523 10999
rect 22756 10996 22784 11036
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 24946 11024 24952 11076
rect 25004 11064 25010 11076
rect 26160 11064 26188 11095
rect 26694 11092 26700 11104
rect 26752 11092 26758 11144
rect 26896 11141 26924 11172
rect 27246 11160 27252 11172
rect 27304 11160 27310 11212
rect 28077 11203 28135 11209
rect 28077 11169 28089 11203
rect 28123 11200 28135 11203
rect 29362 11200 29368 11212
rect 28123 11172 29368 11200
rect 28123 11169 28135 11172
rect 28077 11163 28135 11169
rect 29362 11160 29368 11172
rect 29420 11160 29426 11212
rect 31662 11160 31668 11212
rect 31720 11200 31726 11212
rect 31941 11203 31999 11209
rect 31941 11200 31953 11203
rect 31720 11172 31953 11200
rect 31720 11160 31726 11172
rect 31941 11169 31953 11172
rect 31987 11200 31999 11203
rect 32401 11203 32459 11209
rect 32401 11200 32413 11203
rect 31987 11172 32413 11200
rect 31987 11169 31999 11172
rect 31941 11163 31999 11169
rect 32401 11169 32413 11172
rect 32447 11169 32459 11203
rect 32674 11200 32680 11212
rect 32635 11172 32680 11200
rect 32401 11163 32459 11169
rect 32674 11160 32680 11172
rect 32732 11160 32738 11212
rect 35434 11160 35440 11212
rect 35492 11200 35498 11212
rect 36265 11203 36323 11209
rect 36265 11200 36277 11203
rect 35492 11172 36277 11200
rect 35492 11160 35498 11172
rect 36265 11169 36277 11172
rect 36311 11169 36323 11203
rect 36265 11163 36323 11169
rect 26881 11135 26939 11141
rect 26881 11101 26893 11135
rect 26927 11101 26939 11135
rect 26881 11095 26939 11101
rect 27062 11092 27068 11144
rect 27120 11132 27126 11144
rect 27433 11135 27491 11141
rect 27433 11132 27445 11135
rect 27120 11104 27445 11132
rect 27120 11092 27126 11104
rect 27433 11101 27445 11104
rect 27479 11101 27491 11135
rect 27433 11095 27491 11101
rect 27798 11092 27804 11144
rect 27856 11132 27862 11144
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 27856 11104 28365 11132
rect 27856 11092 27862 11104
rect 28353 11101 28365 11104
rect 28399 11101 28411 11135
rect 28353 11095 28411 11101
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11132 29791 11135
rect 30374 11132 30380 11144
rect 29779 11104 30380 11132
rect 29779 11101 29791 11104
rect 29733 11095 29791 11101
rect 30374 11092 30380 11104
rect 30432 11092 30438 11144
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11132 35035 11135
rect 35805 11135 35863 11141
rect 35805 11132 35817 11135
rect 35023 11104 35817 11132
rect 35023 11101 35035 11104
rect 34977 11095 35035 11101
rect 35805 11101 35817 11104
rect 35851 11132 35863 11135
rect 36078 11132 36084 11144
rect 35851 11104 36084 11132
rect 35851 11101 35863 11104
rect 35805 11095 35863 11101
rect 36078 11092 36084 11104
rect 36136 11092 36142 11144
rect 27816 11064 27844 11092
rect 25004 11036 26188 11064
rect 26252 11036 27844 11064
rect 25004 11024 25010 11036
rect 23382 10996 23388 11008
rect 22756 10968 23388 10996
rect 22465 10959 22523 10965
rect 23382 10956 23388 10968
rect 23440 10956 23446 11008
rect 23658 10956 23664 11008
rect 23716 10996 23722 11008
rect 23753 10999 23811 11005
rect 23753 10996 23765 10999
rect 23716 10968 23765 10996
rect 23716 10956 23722 10968
rect 23753 10965 23765 10968
rect 23799 10965 23811 10999
rect 23753 10959 23811 10965
rect 24302 10956 24308 11008
rect 24360 10996 24366 11008
rect 25406 10996 25412 11008
rect 24360 10968 25412 10996
rect 24360 10956 24366 10968
rect 25406 10956 25412 10968
rect 25464 10996 25470 11008
rect 26252 10996 26280 11036
rect 30926 11024 30932 11076
rect 30984 11024 30990 11076
rect 31570 11024 31576 11076
rect 31628 11064 31634 11076
rect 31665 11067 31723 11073
rect 31665 11064 31677 11067
rect 31628 11036 31677 11064
rect 31628 11024 31634 11036
rect 31665 11033 31677 11036
rect 31711 11033 31723 11067
rect 35618 11064 35624 11076
rect 33902 11036 35624 11064
rect 31665 11027 31723 11033
rect 35618 11024 35624 11036
rect 35676 11024 35682 11076
rect 36449 11067 36507 11073
rect 36449 11033 36461 11067
rect 36495 11064 36507 11067
rect 36630 11064 36636 11076
rect 36495 11036 36636 11064
rect 36495 11033 36507 11036
rect 36449 11027 36507 11033
rect 36630 11024 36636 11036
rect 36688 11024 36694 11076
rect 38105 11067 38163 11073
rect 38105 11033 38117 11067
rect 38151 11064 38163 11067
rect 38194 11064 38200 11076
rect 38151 11036 38200 11064
rect 38151 11033 38163 11036
rect 38105 11027 38163 11033
rect 38194 11024 38200 11036
rect 38252 11024 38258 11076
rect 25464 10968 26280 10996
rect 25464 10956 25470 10968
rect 27246 10956 27252 11008
rect 27304 10996 27310 11008
rect 27890 10996 27896 11008
rect 27304 10968 27896 10996
rect 27304 10956 27310 10968
rect 27890 10956 27896 10968
rect 27948 10996 27954 11008
rect 31018 10996 31024 11008
rect 27948 10968 31024 10996
rect 27948 10956 27954 10968
rect 31018 10956 31024 10968
rect 31076 10956 31082 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 14093 10795 14151 10801
rect 14093 10761 14105 10795
rect 14139 10792 14151 10795
rect 14274 10792 14280 10804
rect 14139 10764 14280 10792
rect 14139 10761 14151 10764
rect 14093 10755 14151 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 15286 10792 15292 10804
rect 14967 10764 15292 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 16448 10764 17233 10792
rect 16448 10752 16454 10764
rect 17221 10761 17233 10764
rect 17267 10761 17279 10795
rect 17221 10755 17279 10761
rect 17957 10795 18015 10801
rect 17957 10761 17969 10795
rect 18003 10792 18015 10795
rect 18046 10792 18052 10804
rect 18003 10764 18052 10792
rect 18003 10761 18015 10764
rect 17957 10755 18015 10761
rect 18046 10752 18052 10764
rect 18104 10792 18110 10804
rect 18325 10795 18383 10801
rect 18104 10764 18276 10792
rect 18104 10752 18110 10764
rect 17126 10724 17132 10736
rect 17087 10696 17132 10724
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 17770 10724 17776 10736
rect 17731 10696 17776 10724
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 18138 10724 18144 10736
rect 18099 10696 18144 10724
rect 18138 10684 18144 10696
rect 18196 10684 18202 10736
rect 18248 10724 18276 10764
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18690 10792 18696 10804
rect 18371 10764 18696 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 21269 10795 21327 10801
rect 21269 10761 21281 10795
rect 21315 10792 21327 10795
rect 22278 10792 22284 10804
rect 21315 10764 22284 10792
rect 21315 10761 21327 10764
rect 21269 10755 21327 10761
rect 19628 10724 19656 10755
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 22557 10795 22615 10801
rect 22557 10761 22569 10795
rect 22603 10792 22615 10795
rect 22738 10792 22744 10804
rect 22603 10764 22744 10792
rect 22603 10761 22615 10764
rect 22557 10755 22615 10761
rect 22738 10752 22744 10764
rect 22796 10752 22802 10804
rect 24489 10795 24547 10801
rect 24136 10764 24440 10792
rect 24136 10736 24164 10764
rect 18248 10696 19656 10724
rect 22649 10727 22707 10733
rect 22649 10693 22661 10727
rect 22695 10724 22707 10727
rect 23198 10724 23204 10736
rect 22695 10696 23204 10724
rect 22695 10693 22707 10696
rect 22649 10687 22707 10693
rect 23198 10684 23204 10696
rect 23256 10684 23262 10736
rect 23934 10724 23940 10736
rect 23308 10696 23940 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14231 10628 14841 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14829 10625 14841 10628
rect 14875 10656 14887 10659
rect 15194 10656 15200 10668
rect 14875 10628 15200 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15436 10628 15761 10656
rect 15436 10616 15442 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16666 10656 16672 10668
rect 15979 10628 16672 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 18104 10628 18149 10656
rect 18248 10628 18981 10656
rect 18104 10616 18110 10628
rect 15654 10588 15660 10600
rect 15615 10560 15660 10588
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 15896 10560 15941 10588
rect 15896 10548 15902 10560
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 18248 10588 18276 10628
rect 18969 10625 18981 10628
rect 19015 10625 19027 10659
rect 19150 10656 19156 10668
rect 19111 10628 19156 10656
rect 18969 10619 19027 10625
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10625 19855 10659
rect 20806 10656 20812 10668
rect 20767 10628 20812 10656
rect 19797 10619 19855 10625
rect 19812 10588 19840 10619
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 21085 10659 21143 10665
rect 21085 10625 21097 10659
rect 21131 10656 21143 10659
rect 22094 10656 22100 10668
rect 21131 10628 22100 10656
rect 21131 10625 21143 10628
rect 21085 10619 21143 10625
rect 22094 10616 22100 10628
rect 22152 10616 22158 10668
rect 22741 10659 22799 10665
rect 22741 10625 22753 10659
rect 22787 10656 22799 10659
rect 23308 10656 23336 10696
rect 23934 10684 23940 10696
rect 23992 10684 23998 10736
rect 24118 10724 24124 10736
rect 24079 10696 24124 10724
rect 24118 10684 24124 10696
rect 24176 10684 24182 10736
rect 24302 10684 24308 10736
rect 24360 10733 24366 10736
rect 24360 10727 24379 10733
rect 24367 10693 24379 10727
rect 24412 10724 24440 10764
rect 24489 10761 24501 10795
rect 24535 10792 24547 10795
rect 25958 10792 25964 10804
rect 24535 10764 25964 10792
rect 24535 10761 24547 10764
rect 24489 10755 24547 10761
rect 25958 10752 25964 10764
rect 26016 10752 26022 10804
rect 27341 10795 27399 10801
rect 27341 10761 27353 10795
rect 27387 10792 27399 10795
rect 27614 10792 27620 10804
rect 27387 10764 27620 10792
rect 27387 10761 27399 10764
rect 27341 10755 27399 10761
rect 27614 10752 27620 10764
rect 27672 10752 27678 10804
rect 29178 10792 29184 10804
rect 29139 10764 29184 10792
rect 29178 10752 29184 10764
rect 29236 10752 29242 10804
rect 30374 10752 30380 10804
rect 30432 10792 30438 10804
rect 30561 10795 30619 10801
rect 30561 10792 30573 10795
rect 30432 10764 30573 10792
rect 30432 10752 30438 10764
rect 30561 10761 30573 10764
rect 30607 10761 30619 10795
rect 31662 10792 31668 10804
rect 30561 10755 30619 10761
rect 31128 10764 31668 10792
rect 25133 10727 25191 10733
rect 25133 10724 25145 10727
rect 24412 10696 25145 10724
rect 24360 10687 24379 10693
rect 25133 10693 25145 10696
rect 25179 10693 25191 10727
rect 25133 10687 25191 10693
rect 25317 10727 25375 10733
rect 25317 10693 25329 10727
rect 25363 10724 25375 10727
rect 25406 10724 25412 10736
rect 25363 10696 25412 10724
rect 25363 10693 25375 10696
rect 25317 10687 25375 10693
rect 24360 10684 24366 10687
rect 25406 10684 25412 10696
rect 25464 10684 25470 10736
rect 26145 10727 26203 10733
rect 26145 10693 26157 10727
rect 26191 10724 26203 10727
rect 26970 10724 26976 10736
rect 26191 10696 26976 10724
rect 26191 10693 26203 10696
rect 26145 10687 26203 10693
rect 26970 10684 26976 10696
rect 27028 10684 27034 10736
rect 28166 10724 28172 10736
rect 27080 10696 28172 10724
rect 22787 10628 23336 10656
rect 22787 10625 22799 10628
rect 22741 10619 22799 10625
rect 23382 10616 23388 10668
rect 23440 10656 23446 10668
rect 23569 10659 23627 10665
rect 23440 10628 23485 10656
rect 23440 10616 23446 10628
rect 23569 10625 23581 10659
rect 23615 10656 23627 10659
rect 23658 10656 23664 10668
rect 23615 10628 23664 10656
rect 23615 10625 23627 10628
rect 23569 10619 23627 10625
rect 23658 10616 23664 10628
rect 23716 10656 23722 10668
rect 24578 10656 24584 10668
rect 23716 10628 24584 10656
rect 23716 10616 23722 10628
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 25222 10656 25228 10668
rect 25135 10628 25228 10656
rect 25222 10616 25228 10628
rect 25280 10656 25286 10668
rect 25590 10656 25596 10668
rect 25280 10628 25596 10656
rect 25280 10616 25286 10628
rect 25590 10616 25596 10628
rect 25648 10656 25654 10668
rect 27080 10656 27108 10696
rect 28166 10684 28172 10696
rect 28224 10684 28230 10736
rect 29270 10684 29276 10736
rect 29328 10724 29334 10736
rect 29822 10724 29828 10736
rect 29328 10696 29828 10724
rect 29328 10684 29334 10696
rect 29822 10684 29828 10696
rect 29880 10724 29886 10736
rect 29880 10696 30420 10724
rect 29880 10684 29886 10696
rect 27246 10656 27252 10668
rect 25648 10628 27108 10656
rect 27207 10628 27252 10656
rect 25648 10616 25654 10628
rect 27246 10616 27252 10628
rect 27304 10616 27310 10668
rect 28074 10616 28080 10668
rect 28132 10656 28138 10668
rect 28132 10628 28580 10656
rect 28132 10616 28138 10628
rect 19886 10588 19892 10600
rect 17736 10560 18276 10588
rect 18984 10560 19892 10588
rect 17736 10548 17742 10560
rect 16850 10480 16856 10532
rect 16908 10520 16914 10532
rect 18984 10520 19012 10560
rect 19886 10548 19892 10560
rect 19944 10588 19950 10600
rect 20622 10588 20628 10600
rect 19944 10560 20628 10588
rect 19944 10548 19950 10560
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 20990 10588 20996 10600
rect 20951 10560 20996 10588
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 22002 10548 22008 10600
rect 22060 10588 22066 10600
rect 23477 10591 23535 10597
rect 23477 10588 23489 10591
rect 22060 10560 23489 10588
rect 22060 10548 22066 10560
rect 23477 10557 23489 10560
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 24670 10548 24676 10600
rect 24728 10588 24734 10600
rect 24728 10560 26280 10588
rect 24728 10548 24734 10560
rect 16908 10492 19012 10520
rect 19061 10523 19119 10529
rect 16908 10480 16914 10492
rect 19061 10489 19073 10523
rect 19107 10520 19119 10523
rect 19107 10492 20852 10520
rect 19107 10489 19119 10492
rect 19061 10483 19119 10489
rect 15473 10455 15531 10461
rect 15473 10421 15485 10455
rect 15519 10452 15531 10455
rect 15562 10452 15568 10464
rect 15519 10424 15568 10452
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16758 10412 16764 10464
rect 16816 10452 16822 10464
rect 19426 10452 19432 10464
rect 16816 10424 19432 10452
rect 16816 10412 16822 10424
rect 19426 10412 19432 10424
rect 19484 10452 19490 10464
rect 19702 10452 19708 10464
rect 19484 10424 19708 10452
rect 19484 10412 19490 10424
rect 19702 10412 19708 10424
rect 19760 10452 19766 10464
rect 20530 10452 20536 10464
rect 19760 10424 20536 10452
rect 19760 10412 19766 10424
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 20824 10461 20852 10492
rect 20898 10480 20904 10532
rect 20956 10520 20962 10532
rect 22373 10523 22431 10529
rect 22373 10520 22385 10523
rect 20956 10492 22385 10520
rect 20956 10480 20962 10492
rect 22373 10489 22385 10492
rect 22419 10489 22431 10523
rect 22373 10483 22431 10489
rect 23382 10480 23388 10532
rect 23440 10520 23446 10532
rect 24118 10520 24124 10532
rect 23440 10492 24124 10520
rect 23440 10480 23446 10492
rect 24118 10480 24124 10492
rect 24176 10520 24182 10532
rect 24946 10520 24952 10532
rect 24176 10492 24952 10520
rect 24176 10480 24182 10492
rect 24946 10480 24952 10492
rect 25004 10480 25010 10532
rect 25501 10523 25559 10529
rect 25501 10489 25513 10523
rect 25547 10520 25559 10523
rect 26142 10520 26148 10532
rect 25547 10492 26148 10520
rect 25547 10489 25559 10492
rect 25501 10483 25559 10489
rect 26142 10480 26148 10492
rect 26200 10480 26206 10532
rect 26252 10520 26280 10560
rect 28166 10548 28172 10600
rect 28224 10588 28230 10600
rect 28445 10591 28503 10597
rect 28445 10588 28457 10591
rect 28224 10560 28457 10588
rect 28224 10548 28230 10560
rect 28445 10557 28457 10560
rect 28491 10557 28503 10591
rect 28552 10588 28580 10628
rect 28626 10616 28632 10668
rect 28684 10656 28690 10668
rect 30392 10665 30420 10696
rect 30834 10684 30840 10736
rect 30892 10724 30898 10736
rect 31128 10733 31156 10764
rect 31662 10752 31668 10764
rect 31720 10792 31726 10804
rect 33870 10792 33876 10804
rect 31720 10752 31754 10792
rect 33831 10764 33876 10792
rect 33870 10752 33876 10764
rect 33928 10752 33934 10804
rect 31113 10727 31171 10733
rect 31113 10724 31125 10727
rect 30892 10696 31125 10724
rect 30892 10684 30898 10696
rect 31113 10693 31125 10696
rect 31159 10693 31171 10727
rect 31113 10687 31171 10693
rect 31297 10727 31355 10733
rect 31297 10693 31309 10727
rect 31343 10724 31355 10727
rect 31386 10724 31392 10736
rect 31343 10696 31392 10724
rect 31343 10693 31355 10696
rect 31297 10687 31355 10693
rect 31386 10684 31392 10696
rect 31444 10684 31450 10736
rect 31726 10724 31754 10752
rect 31726 10696 32168 10724
rect 32140 10665 32168 10696
rect 33410 10684 33416 10736
rect 33468 10684 33474 10736
rect 36538 10724 36544 10736
rect 36499 10696 36544 10724
rect 36538 10684 36544 10696
rect 36596 10684 36602 10736
rect 28721 10659 28779 10665
rect 28721 10656 28733 10659
rect 28684 10628 28733 10656
rect 28684 10616 28690 10628
rect 28721 10625 28733 10628
rect 28767 10656 28779 10659
rect 29365 10659 29423 10665
rect 29365 10656 29377 10659
rect 28767 10628 29377 10656
rect 28767 10625 28779 10628
rect 28721 10619 28779 10625
rect 29365 10625 29377 10628
rect 29411 10625 29423 10659
rect 29365 10619 29423 10625
rect 29733 10659 29791 10665
rect 29733 10625 29745 10659
rect 29779 10625 29791 10659
rect 29733 10619 29791 10625
rect 30377 10659 30435 10665
rect 30377 10625 30389 10659
rect 30423 10625 30435 10659
rect 30377 10619 30435 10625
rect 32125 10659 32183 10665
rect 32125 10625 32137 10659
rect 32171 10625 32183 10659
rect 32125 10619 32183 10625
rect 37369 10659 37427 10665
rect 37369 10625 37381 10659
rect 37415 10656 37427 10659
rect 38562 10656 38568 10668
rect 37415 10628 38568 10656
rect 37415 10625 37427 10628
rect 37369 10619 37427 10625
rect 29748 10588 29776 10619
rect 38562 10616 38568 10628
rect 38620 10616 38626 10668
rect 28552 10560 29776 10588
rect 29825 10591 29883 10597
rect 28445 10551 28503 10557
rect 29825 10557 29837 10591
rect 29871 10588 29883 10591
rect 30190 10588 30196 10600
rect 29871 10560 30196 10588
rect 29871 10557 29883 10560
rect 29825 10551 29883 10557
rect 30190 10548 30196 10560
rect 30248 10548 30254 10600
rect 31662 10548 31668 10600
rect 31720 10588 31726 10600
rect 32401 10591 32459 10597
rect 32401 10588 32413 10591
rect 31720 10560 32413 10588
rect 31720 10548 31726 10560
rect 32401 10557 32413 10560
rect 32447 10557 32459 10591
rect 35802 10588 35808 10600
rect 35763 10560 35808 10588
rect 32401 10551 32459 10557
rect 35802 10548 35808 10560
rect 35860 10548 35866 10600
rect 36722 10588 36728 10600
rect 36683 10560 36728 10588
rect 36722 10548 36728 10560
rect 36780 10548 36786 10600
rect 32122 10520 32128 10532
rect 26252 10492 32128 10520
rect 32122 10480 32128 10492
rect 32180 10480 32186 10532
rect 20809 10455 20867 10461
rect 20809 10421 20821 10455
rect 20855 10452 20867 10455
rect 21542 10452 21548 10464
rect 20855 10424 21548 10452
rect 20855 10421 20867 10424
rect 20809 10415 20867 10421
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 22738 10412 22744 10464
rect 22796 10452 22802 10464
rect 22925 10455 22983 10461
rect 22925 10452 22937 10455
rect 22796 10424 22937 10452
rect 22796 10412 22802 10424
rect 22925 10421 22937 10424
rect 22971 10421 22983 10455
rect 22925 10415 22983 10421
rect 24305 10455 24363 10461
rect 24305 10421 24317 10455
rect 24351 10452 24363 10455
rect 25222 10452 25228 10464
rect 24351 10424 25228 10452
rect 24351 10421 24363 10424
rect 24305 10415 24363 10421
rect 25222 10412 25228 10424
rect 25280 10412 25286 10464
rect 26053 10455 26111 10461
rect 26053 10421 26065 10455
rect 26099 10452 26111 10455
rect 26234 10452 26240 10464
rect 26099 10424 26240 10452
rect 26099 10421 26111 10424
rect 26053 10415 26111 10421
rect 26234 10412 26240 10424
rect 26292 10412 26298 10464
rect 29362 10452 29368 10464
rect 29323 10424 29368 10452
rect 29362 10412 29368 10424
rect 29420 10412 29426 10464
rect 36446 10412 36452 10464
rect 36504 10452 36510 10464
rect 37461 10455 37519 10461
rect 37461 10452 37473 10455
rect 36504 10424 37473 10452
rect 36504 10412 36510 10424
rect 37461 10421 37473 10424
rect 37507 10421 37519 10455
rect 37461 10415 37519 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 17313 10251 17371 10257
rect 17313 10217 17325 10251
rect 17359 10248 17371 10251
rect 17586 10248 17592 10260
rect 17359 10220 17592 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 17586 10208 17592 10220
rect 17644 10248 17650 10260
rect 17644 10220 18000 10248
rect 17644 10208 17650 10220
rect 16850 10140 16856 10192
rect 16908 10140 16914 10192
rect 16868 10112 16896 10140
rect 17972 10121 18000 10220
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 18104 10220 18337 10248
rect 18104 10208 18110 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 19702 10248 19708 10260
rect 19663 10220 19708 10248
rect 18325 10211 18383 10217
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 19978 10248 19984 10260
rect 19939 10220 19984 10248
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20530 10248 20536 10260
rect 20491 10220 20536 10248
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 20990 10208 20996 10260
rect 21048 10248 21054 10260
rect 21085 10251 21143 10257
rect 21085 10248 21097 10251
rect 21048 10220 21097 10248
rect 21048 10208 21054 10220
rect 21085 10217 21097 10220
rect 21131 10217 21143 10251
rect 21085 10211 21143 10217
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 22704 10220 22937 10248
rect 22704 10208 22710 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 23566 10248 23572 10260
rect 23527 10220 23572 10248
rect 22925 10211 22983 10217
rect 23566 10208 23572 10220
rect 23624 10208 23630 10260
rect 27525 10251 27583 10257
rect 27525 10248 27537 10251
rect 23860 10220 27537 10248
rect 20070 10180 20076 10192
rect 18064 10152 20076 10180
rect 17957 10115 18015 10121
rect 16868 10084 16988 10112
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14921 10047 14979 10053
rect 14921 10044 14933 10047
rect 14139 10016 14933 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 14921 10013 14933 10016
rect 14967 10044 14979 10047
rect 15194 10044 15200 10056
rect 14967 10016 15200 10044
rect 14967 10013 14979 10016
rect 14921 10007 14979 10013
rect 15194 10004 15200 10016
rect 15252 10004 15258 10056
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 16025 10047 16083 10053
rect 16025 10044 16037 10047
rect 15436 10016 16037 10044
rect 15436 10004 15442 10016
rect 16025 10013 16037 10016
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10044 16359 10047
rect 16574 10044 16580 10056
rect 16347 10016 16580 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 16040 9976 16068 10007
rect 16574 10004 16580 10016
rect 16632 10044 16638 10056
rect 16960 10053 16988 10084
rect 17957 10081 17969 10115
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16632 10016 16865 10044
rect 16632 10004 16638 10016
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 17310 10044 17316 10056
rect 17271 10016 17316 10044
rect 16945 10007 17003 10013
rect 17310 10004 17316 10016
rect 17368 10044 17374 10056
rect 18064 10044 18092 10152
rect 20070 10140 20076 10152
rect 20128 10140 20134 10192
rect 22094 10140 22100 10192
rect 22152 10180 22158 10192
rect 22189 10183 22247 10189
rect 22189 10180 22201 10183
rect 22152 10152 22201 10180
rect 22152 10140 22158 10152
rect 22189 10149 22201 10152
rect 22235 10149 22247 10183
rect 22189 10143 22247 10149
rect 18782 10072 18788 10124
rect 18840 10112 18846 10124
rect 20809 10115 20867 10121
rect 18840 10084 19840 10112
rect 18840 10072 18846 10084
rect 17368 10016 18092 10044
rect 18141 10047 18199 10053
rect 17368 10004 17374 10016
rect 18141 10013 18153 10047
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18156 9976 18184 10007
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 19812 10053 19840 10084
rect 20809 10081 20821 10115
rect 20855 10112 20867 10115
rect 22002 10112 22008 10124
rect 20855 10084 22008 10112
rect 20855 10081 20867 10084
rect 20809 10075 20867 10081
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 22738 10112 22744 10124
rect 22699 10084 22744 10112
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 19024 10016 19349 10044
rect 19024 10004 19030 10016
rect 19337 10013 19349 10016
rect 19383 10013 19395 10047
rect 19337 10007 19395 10013
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10044 19855 10047
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 19843 10016 20913 10044
rect 19843 10013 19855 10016
rect 19797 10007 19855 10013
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 18322 9976 18328 9988
rect 16040 9948 18328 9976
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 18874 9936 18880 9988
rect 18932 9976 18938 9988
rect 19150 9976 19156 9988
rect 18932 9948 19156 9976
rect 18932 9936 18938 9948
rect 19150 9936 19156 9948
rect 19208 9976 19214 9988
rect 19444 9976 19472 10007
rect 23474 10004 23480 10056
rect 23532 10044 23538 10056
rect 23860 10053 23888 10220
rect 27525 10217 27537 10220
rect 27571 10217 27583 10251
rect 27798 10248 27804 10260
rect 27759 10220 27804 10248
rect 27525 10211 27583 10217
rect 27798 10208 27804 10220
rect 27856 10208 27862 10260
rect 27890 10208 27896 10260
rect 27948 10248 27954 10260
rect 30190 10248 30196 10260
rect 27948 10220 30196 10248
rect 27948 10208 27954 10220
rect 30190 10208 30196 10220
rect 30248 10208 30254 10260
rect 30926 10248 30932 10260
rect 30887 10220 30932 10248
rect 30926 10208 30932 10220
rect 30984 10208 30990 10260
rect 31662 10248 31668 10260
rect 31623 10220 31668 10248
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 32122 10208 32128 10260
rect 32180 10248 32186 10260
rect 32217 10251 32275 10257
rect 32217 10248 32229 10251
rect 32180 10220 32229 10248
rect 32180 10208 32186 10220
rect 32217 10217 32229 10220
rect 32263 10217 32275 10251
rect 32217 10211 32275 10217
rect 34977 10251 35035 10257
rect 34977 10217 34989 10251
rect 35023 10248 35035 10251
rect 35342 10248 35348 10260
rect 35023 10220 35348 10248
rect 35023 10217 35035 10220
rect 34977 10211 35035 10217
rect 35342 10208 35348 10220
rect 35400 10208 35406 10260
rect 35618 10248 35624 10260
rect 35579 10220 35624 10248
rect 35618 10208 35624 10220
rect 35676 10208 35682 10260
rect 26326 10140 26332 10192
rect 26384 10180 26390 10192
rect 28994 10180 29000 10192
rect 26384 10152 29000 10180
rect 26384 10140 26390 10152
rect 28994 10140 29000 10152
rect 29052 10140 29058 10192
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10112 25007 10115
rect 26234 10112 26240 10124
rect 24995 10084 26240 10112
rect 24995 10081 25007 10084
rect 24949 10075 25007 10081
rect 26234 10072 26240 10084
rect 26292 10112 26298 10124
rect 27522 10112 27528 10124
rect 26292 10084 27528 10112
rect 26292 10072 26298 10084
rect 27522 10072 27528 10084
rect 27580 10072 27586 10124
rect 28166 10112 28172 10124
rect 28127 10084 28172 10112
rect 28166 10072 28172 10084
rect 28224 10072 28230 10124
rect 34149 10115 34207 10121
rect 30852 10084 32996 10112
rect 23569 10047 23627 10053
rect 23569 10044 23581 10047
rect 23532 10016 23581 10044
rect 23532 10004 23538 10016
rect 23569 10013 23581 10016
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10013 23903 10047
rect 23845 10007 23903 10013
rect 27709 10047 27767 10053
rect 27709 10013 27721 10047
rect 27755 10044 27767 10047
rect 27890 10044 27896 10056
rect 27755 10016 27896 10044
rect 27755 10013 27767 10016
rect 27709 10007 27767 10013
rect 20438 9976 20444 9988
rect 19208 9948 19472 9976
rect 20399 9948 20444 9976
rect 19208 9936 19214 9948
rect 20438 9936 20444 9948
rect 20496 9936 20502 9988
rect 22186 9976 22192 9988
rect 22147 9948 22192 9976
rect 22186 9936 22192 9948
rect 22244 9936 22250 9988
rect 23676 9976 23704 10007
rect 27890 10004 27896 10016
rect 27948 10004 27954 10056
rect 28074 10044 28080 10056
rect 28035 10016 28080 10044
rect 28074 10004 28080 10016
rect 28132 10004 28138 10056
rect 28258 10004 28264 10056
rect 28316 10044 28322 10056
rect 28721 10047 28779 10053
rect 28721 10044 28733 10047
rect 28316 10016 28733 10044
rect 28316 10004 28322 10016
rect 28721 10013 28733 10016
rect 28767 10013 28779 10047
rect 28721 10007 28779 10013
rect 28813 10047 28871 10053
rect 28813 10013 28825 10047
rect 28859 10044 28871 10047
rect 29638 10044 29644 10056
rect 28859 10016 29644 10044
rect 28859 10013 28871 10016
rect 28813 10007 28871 10013
rect 29638 10004 29644 10016
rect 29696 10004 29702 10056
rect 29822 10044 29828 10056
rect 29783 10016 29828 10044
rect 29822 10004 29828 10016
rect 29880 10004 29886 10056
rect 30374 10004 30380 10056
rect 30432 10044 30438 10056
rect 30852 10053 30880 10084
rect 32968 10056 32996 10084
rect 34149 10081 34161 10115
rect 34195 10112 34207 10115
rect 36265 10115 36323 10121
rect 36265 10112 36277 10115
rect 34195 10084 36277 10112
rect 34195 10081 34207 10084
rect 34149 10075 34207 10081
rect 36265 10081 36277 10084
rect 36311 10081 36323 10115
rect 36446 10112 36452 10124
rect 36407 10084 36452 10112
rect 36265 10075 36323 10081
rect 36446 10072 36452 10084
rect 36504 10072 36510 10124
rect 38102 10112 38108 10124
rect 38063 10084 38108 10112
rect 38102 10072 38108 10084
rect 38160 10072 38166 10124
rect 30837 10047 30895 10053
rect 30837 10044 30849 10047
rect 30432 10016 30849 10044
rect 30432 10004 30438 10016
rect 30837 10013 30849 10016
rect 30883 10013 30895 10047
rect 30837 10007 30895 10013
rect 31481 10047 31539 10053
rect 31481 10013 31493 10047
rect 31527 10044 31539 10047
rect 31754 10044 31760 10056
rect 31527 10016 31760 10044
rect 31527 10013 31539 10016
rect 31481 10007 31539 10013
rect 31754 10004 31760 10016
rect 31812 10004 31818 10056
rect 32125 10047 32183 10053
rect 32125 10013 32137 10047
rect 32171 10013 32183 10047
rect 32125 10007 32183 10013
rect 25222 9976 25228 9988
rect 23676 9948 23888 9976
rect 25183 9948 25228 9976
rect 23860 9920 23888 9948
rect 25222 9936 25228 9948
rect 25280 9936 25286 9988
rect 28534 9976 28540 9988
rect 26450 9948 28540 9976
rect 28534 9936 28540 9948
rect 28592 9936 28598 9988
rect 28994 9936 29000 9988
rect 29052 9976 29058 9988
rect 29052 9948 29097 9976
rect 29052 9936 29058 9948
rect 31018 9936 31024 9988
rect 31076 9976 31082 9988
rect 32140 9976 32168 10007
rect 32950 10004 32956 10056
rect 33008 10044 33014 10056
rect 34885 10047 34943 10053
rect 34885 10044 34897 10047
rect 33008 10016 34897 10044
rect 33008 10004 33014 10016
rect 34885 10013 34897 10016
rect 34931 10044 34943 10047
rect 35529 10047 35587 10053
rect 35529 10044 35541 10047
rect 34931 10016 35541 10044
rect 34931 10013 34943 10016
rect 34885 10007 34943 10013
rect 35529 10013 35541 10016
rect 35575 10013 35587 10047
rect 35529 10007 35587 10013
rect 31076 9948 32168 9976
rect 31076 9936 31082 9948
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 14185 9911 14243 9917
rect 14185 9908 14197 9911
rect 14148 9880 14197 9908
rect 14148 9868 14154 9880
rect 14185 9877 14197 9880
rect 14231 9877 14243 9911
rect 14826 9908 14832 9920
rect 14787 9880 14832 9908
rect 14185 9871 14243 9877
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 17497 9911 17555 9917
rect 17497 9877 17509 9911
rect 17543 9908 17555 9911
rect 19242 9908 19248 9920
rect 17543 9880 19248 9908
rect 17543 9877 17555 9880
rect 17497 9871 17555 9877
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 22646 9908 22652 9920
rect 22607 9880 22652 9908
rect 22646 9868 22652 9880
rect 22704 9868 22710 9920
rect 23382 9908 23388 9920
rect 23343 9880 23388 9908
rect 23382 9868 23388 9880
rect 23440 9868 23446 9920
rect 23842 9868 23848 9920
rect 23900 9868 23906 9920
rect 26694 9908 26700 9920
rect 26655 9880 26700 9908
rect 26694 9868 26700 9880
rect 26752 9868 26758 9920
rect 27890 9868 27896 9920
rect 27948 9908 27954 9920
rect 28721 9911 28779 9917
rect 28721 9908 28733 9911
rect 27948 9880 28733 9908
rect 27948 9868 27954 9880
rect 28721 9877 28733 9880
rect 28767 9877 28779 9911
rect 28721 9871 28779 9877
rect 29641 9911 29699 9917
rect 29641 9877 29653 9911
rect 29687 9908 29699 9911
rect 30374 9908 30380 9920
rect 29687 9880 30380 9908
rect 29687 9877 29699 9880
rect 29641 9871 29699 9877
rect 30374 9868 30380 9880
rect 30432 9868 30438 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 18046 9704 18052 9716
rect 18007 9676 18052 9704
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 18230 9704 18236 9716
rect 18191 9676 18236 9704
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 19061 9707 19119 9713
rect 19061 9673 19073 9707
rect 19107 9673 19119 9707
rect 20806 9704 20812 9716
rect 20767 9676 20812 9704
rect 19061 9667 19119 9673
rect 14090 9596 14096 9648
rect 14148 9596 14154 9648
rect 16850 9636 16856 9648
rect 15856 9608 16856 9636
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 15856 9577 15884 9608
rect 16850 9596 16856 9608
rect 16908 9596 16914 9648
rect 16942 9596 16948 9648
rect 17000 9596 17006 9648
rect 17865 9639 17923 9645
rect 17865 9605 17877 9639
rect 17911 9636 17923 9639
rect 17954 9636 17960 9648
rect 17911 9608 17960 9636
rect 17911 9605 17923 9608
rect 17865 9599 17923 9605
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 18141 9639 18199 9645
rect 18141 9605 18153 9639
rect 18187 9636 18199 9639
rect 18690 9636 18696 9648
rect 18187 9608 18696 9636
rect 18187 9605 18199 9608
rect 18141 9599 18199 9605
rect 18690 9596 18696 9608
rect 18748 9596 18754 9648
rect 19076 9636 19104 9667
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 22097 9707 22155 9713
rect 20956 9676 21404 9704
rect 20956 9664 20962 9676
rect 19076 9608 19196 9636
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 15841 9531 15899 9537
rect 16132 9540 16681 9568
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 13446 9500 13452 9512
rect 13403 9472 13452 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 16132 9509 16160 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16960 9568 16988 9596
rect 19168 9580 19196 9608
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 21269 9639 21327 9645
rect 21269 9636 21281 9639
rect 19300 9608 21281 9636
rect 19300 9596 19306 9608
rect 21269 9605 21281 9608
rect 21315 9605 21327 9639
rect 21376 9636 21404 9676
rect 22097 9673 22109 9707
rect 22143 9704 22155 9707
rect 22143 9676 22232 9704
rect 22143 9673 22155 9676
rect 22097 9667 22155 9673
rect 22204 9636 22232 9676
rect 25222 9664 25228 9716
rect 25280 9704 25286 9716
rect 25409 9707 25467 9713
rect 25409 9704 25421 9707
rect 25280 9676 25421 9704
rect 25280 9664 25286 9676
rect 25409 9673 25421 9676
rect 25455 9673 25467 9707
rect 28258 9704 28264 9716
rect 25409 9667 25467 9673
rect 27356 9676 28264 9704
rect 22554 9636 22560 9648
rect 21376 9608 22094 9636
rect 22204 9608 22560 9636
rect 21269 9599 21327 9605
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 16960 9540 17141 9568
rect 16669 9531 16727 9537
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 18874 9568 18880 9580
rect 17460 9540 18880 9568
rect 17460 9528 17466 9540
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 19024 9540 19069 9568
rect 19024 9528 19030 9540
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 19705 9571 19763 9577
rect 19208 9540 19380 9568
rect 19208 9528 19214 9540
rect 16117 9503 16175 9509
rect 16117 9469 16129 9503
rect 16163 9469 16175 9503
rect 16117 9463 16175 9469
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 16132 9432 16160 9463
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16632 9472 16957 9500
rect 16632 9460 16638 9472
rect 16945 9469 16957 9472
rect 16991 9500 17003 9503
rect 17218 9500 17224 9512
rect 16991 9472 17224 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 18104 9472 19257 9500
rect 18104 9460 18110 9472
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19352 9500 19380 9540
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 19886 9568 19892 9580
rect 19751 9540 19892 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20165 9571 20223 9577
rect 20165 9568 20177 9571
rect 20128 9540 20177 9568
rect 20128 9528 20134 9540
rect 20165 9537 20177 9540
rect 20211 9537 20223 9571
rect 20165 9531 20223 9537
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9568 21051 9571
rect 21450 9568 21456 9580
rect 21039 9540 21456 9568
rect 21039 9537 21051 9540
rect 20993 9531 21051 9537
rect 21450 9528 21456 9540
rect 21508 9528 21514 9580
rect 22066 9568 22094 9608
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 22741 9639 22799 9645
rect 22741 9605 22753 9639
rect 22787 9636 22799 9639
rect 23382 9636 23388 9648
rect 22787 9608 23388 9636
rect 22787 9605 22799 9608
rect 22741 9599 22799 9605
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 25682 9636 25688 9648
rect 24044 9608 25688 9636
rect 22462 9568 22468 9580
rect 22066 9540 22468 9568
rect 22462 9528 22468 9540
rect 22520 9528 22526 9580
rect 24044 9577 24072 9608
rect 25682 9596 25688 9608
rect 25740 9596 25746 9648
rect 25958 9596 25964 9648
rect 26016 9636 26022 9648
rect 27356 9636 27384 9676
rect 28258 9664 28264 9676
rect 28316 9664 28322 9716
rect 30190 9664 30196 9716
rect 30248 9704 30254 9716
rect 30377 9707 30435 9713
rect 30377 9704 30389 9707
rect 30248 9676 30389 9704
rect 30248 9664 30254 9676
rect 30377 9673 30389 9676
rect 30423 9673 30435 9707
rect 30377 9667 30435 9673
rect 27522 9636 27528 9648
rect 26016 9608 27384 9636
rect 27483 9608 27528 9636
rect 26016 9596 26022 9608
rect 23661 9571 23719 9577
rect 23661 9537 23673 9571
rect 23707 9568 23719 9571
rect 24029 9571 24087 9577
rect 23707 9540 23980 9568
rect 23707 9537 23719 9540
rect 23661 9531 23719 9537
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 19352 9472 19993 9500
rect 19245 9463 19303 9469
rect 19981 9469 19993 9472
rect 20027 9469 20039 9503
rect 20898 9500 20904 9512
rect 19981 9463 20039 9469
rect 20272 9472 20904 9500
rect 15528 9404 16160 9432
rect 18417 9435 18475 9441
rect 15528 9392 15534 9404
rect 18417 9401 18429 9435
rect 18463 9432 18475 9435
rect 18598 9432 18604 9444
rect 18463 9404 18604 9432
rect 18463 9401 18475 9404
rect 18417 9395 18475 9401
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 19153 9435 19211 9441
rect 19153 9401 19165 9435
rect 19199 9432 19211 9435
rect 20272 9432 20300 9472
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 21174 9460 21180 9512
rect 21232 9500 21238 9512
rect 21232 9472 21277 9500
rect 21232 9460 21238 9472
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 22152 9472 22385 9500
rect 22152 9460 22158 9472
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 23474 9460 23480 9512
rect 23532 9460 23538 9512
rect 19199 9404 20300 9432
rect 20349 9435 20407 9441
rect 19199 9401 19211 9404
rect 19153 9395 19211 9401
rect 20349 9401 20361 9435
rect 20395 9432 20407 9435
rect 23492 9432 23520 9460
rect 23750 9432 23756 9444
rect 20395 9404 23520 9432
rect 23584 9404 23756 9432
rect 20395 9401 20407 9404
rect 20349 9395 20407 9401
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1452 9336 1593 9364
rect 1452 9324 1458 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 2869 9367 2927 9373
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 4062 9364 4068 9376
rect 2915 9336 4068 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 16574 9364 16580 9376
rect 14875 9336 16580 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 16758 9364 16764 9376
rect 16719 9336 16764 9364
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 17313 9367 17371 9373
rect 17313 9333 17325 9367
rect 17359 9364 17371 9367
rect 19334 9364 19340 9376
rect 17359 9336 19340 9364
rect 17359 9333 17371 9336
rect 17313 9327 17371 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19978 9364 19984 9376
rect 19939 9336 19984 9364
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 20993 9367 21051 9373
rect 20993 9364 21005 9367
rect 20956 9336 21005 9364
rect 20956 9324 20962 9336
rect 20993 9333 21005 9336
rect 21039 9333 21051 9367
rect 20993 9327 21051 9333
rect 21542 9324 21548 9376
rect 21600 9364 21606 9376
rect 22465 9367 22523 9373
rect 22465 9364 22477 9367
rect 21600 9336 22477 9364
rect 21600 9324 21606 9336
rect 22465 9333 22477 9336
rect 22511 9333 22523 9367
rect 22465 9327 22523 9333
rect 22603 9367 22661 9373
rect 22603 9333 22615 9367
rect 22649 9364 22661 9367
rect 22738 9364 22744 9376
rect 22649 9336 22744 9364
rect 22649 9333 22661 9336
rect 22603 9327 22661 9333
rect 22738 9324 22744 9336
rect 22796 9324 22802 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23584 9364 23612 9404
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 23952 9432 23980 9540
rect 24029 9537 24041 9571
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 24118 9528 24124 9580
rect 24176 9568 24182 9580
rect 25225 9571 25283 9577
rect 24176 9540 24221 9568
rect 24176 9528 24182 9540
rect 25225 9537 25237 9571
rect 25271 9568 25283 9571
rect 25314 9568 25320 9580
rect 25271 9540 25320 9568
rect 25271 9537 25283 9540
rect 25225 9531 25283 9537
rect 25314 9528 25320 9540
rect 25372 9528 25378 9580
rect 25866 9528 25872 9580
rect 25924 9568 25930 9580
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 25924 9540 26065 9568
rect 25924 9528 25930 9540
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26418 9528 26424 9580
rect 26476 9568 26482 9580
rect 27154 9568 27160 9580
rect 26476 9540 27160 9568
rect 26476 9528 26482 9540
rect 27154 9528 27160 9540
rect 27212 9528 27218 9580
rect 27264 9577 27292 9608
rect 27522 9596 27528 9608
rect 27580 9596 27586 9648
rect 27617 9639 27675 9645
rect 27617 9605 27629 9639
rect 27663 9636 27675 9639
rect 27893 9639 27951 9645
rect 27663 9608 27844 9636
rect 27663 9605 27675 9608
rect 27617 9599 27675 9605
rect 27430 9577 27436 9580
rect 27249 9571 27307 9577
rect 27249 9537 27261 9571
rect 27295 9537 27307 9571
rect 27407 9571 27436 9577
rect 27407 9568 27419 9571
rect 27343 9540 27419 9568
rect 27249 9531 27307 9537
rect 27407 9537 27419 9540
rect 27407 9531 27436 9537
rect 27430 9528 27436 9531
rect 27488 9528 27494 9580
rect 27709 9571 27767 9577
rect 27709 9537 27721 9571
rect 27755 9537 27767 9571
rect 27709 9531 27767 9537
rect 24670 9460 24676 9512
rect 24728 9500 24734 9512
rect 24949 9503 25007 9509
rect 24949 9500 24961 9503
rect 24728 9472 24961 9500
rect 24728 9460 24734 9472
rect 24949 9469 24961 9472
rect 24995 9500 25007 9503
rect 25958 9500 25964 9512
rect 24995 9472 25176 9500
rect 25919 9472 25964 9500
rect 24995 9469 25007 9472
rect 24949 9463 25007 9469
rect 24118 9432 24124 9444
rect 23952 9404 24124 9432
rect 24118 9392 24124 9404
rect 24176 9392 24182 9444
rect 23523 9336 23612 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23658 9324 23664 9376
rect 23716 9364 23722 9376
rect 25038 9364 25044 9376
rect 23716 9336 23761 9364
rect 24999 9336 25044 9364
rect 23716 9324 23722 9336
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 25148 9364 25176 9472
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 26142 9500 26148 9512
rect 26103 9472 26148 9500
rect 26142 9460 26148 9472
rect 26200 9460 26206 9512
rect 26234 9460 26240 9512
rect 26292 9500 26298 9512
rect 26292 9472 26337 9500
rect 26292 9460 26298 9472
rect 26510 9460 26516 9512
rect 26568 9500 26574 9512
rect 27448 9500 27476 9528
rect 26568 9472 27476 9500
rect 26568 9460 26574 9472
rect 26421 9435 26479 9441
rect 26421 9401 26433 9435
rect 26467 9432 26479 9435
rect 27724 9432 27752 9531
rect 27816 9500 27844 9608
rect 27893 9605 27905 9639
rect 27939 9636 27951 9639
rect 28905 9639 28963 9645
rect 28905 9636 28917 9639
rect 27939 9608 28917 9636
rect 27939 9605 27951 9608
rect 27893 9599 27951 9605
rect 28905 9605 28917 9608
rect 28951 9605 28963 9639
rect 28905 9599 28963 9605
rect 30466 9596 30472 9648
rect 30524 9636 30530 9648
rect 30929 9639 30987 9645
rect 30929 9636 30941 9639
rect 30524 9608 30941 9636
rect 30524 9596 30530 9608
rect 30929 9605 30941 9608
rect 30975 9605 30987 9639
rect 36630 9636 36636 9648
rect 36591 9608 36636 9636
rect 30929 9599 30987 9605
rect 36630 9596 36636 9608
rect 36688 9596 36694 9648
rect 30006 9528 30012 9580
rect 30064 9528 30070 9580
rect 31018 9568 31024 9580
rect 30979 9540 31024 9568
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 35805 9571 35863 9577
rect 35805 9537 35817 9571
rect 35851 9568 35863 9571
rect 35986 9568 35992 9580
rect 35851 9540 35992 9568
rect 35851 9537 35863 9540
rect 35805 9531 35863 9537
rect 35986 9528 35992 9540
rect 36044 9528 36050 9580
rect 36725 9571 36783 9577
rect 36725 9537 36737 9571
rect 36771 9568 36783 9571
rect 36998 9568 37004 9580
rect 36771 9540 37004 9568
rect 36771 9537 36783 9540
rect 36725 9531 36783 9537
rect 36998 9528 37004 9540
rect 37056 9528 37062 9580
rect 37461 9571 37519 9577
rect 37461 9537 37473 9571
rect 37507 9568 37519 9571
rect 38378 9568 38384 9580
rect 37507 9540 38384 9568
rect 37507 9537 37519 9540
rect 37461 9531 37519 9537
rect 38378 9528 38384 9540
rect 38436 9528 38442 9580
rect 27890 9500 27896 9512
rect 27816 9472 27896 9500
rect 27890 9460 27896 9472
rect 27948 9460 27954 9512
rect 28626 9500 28632 9512
rect 28587 9472 28632 9500
rect 28626 9460 28632 9472
rect 28684 9460 28690 9512
rect 35161 9503 35219 9509
rect 35161 9469 35173 9503
rect 35207 9500 35219 9503
rect 36170 9500 36176 9512
rect 35207 9472 36176 9500
rect 35207 9469 35219 9472
rect 35161 9463 35219 9469
rect 36170 9460 36176 9472
rect 36228 9460 36234 9512
rect 26467 9404 27752 9432
rect 34149 9435 34207 9441
rect 26467 9401 26479 9404
rect 26421 9395 26479 9401
rect 34149 9401 34161 9435
rect 34195 9432 34207 9435
rect 36262 9432 36268 9444
rect 34195 9404 36268 9432
rect 34195 9401 34207 9404
rect 34149 9395 34207 9401
rect 36262 9392 36268 9404
rect 36320 9392 36326 9444
rect 26970 9364 26976 9376
rect 25148 9336 26976 9364
rect 26970 9324 26976 9336
rect 27028 9324 27034 9376
rect 37553 9367 37611 9373
rect 37553 9333 37565 9367
rect 37599 9364 37611 9367
rect 37918 9364 37924 9376
rect 37599 9336 37924 9364
rect 37599 9333 37611 9336
rect 37553 9327 37611 9333
rect 37918 9324 37924 9336
rect 37976 9324 37982 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 13446 9160 13452 9172
rect 13407 9132 13452 9160
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 15470 9160 15476 9172
rect 14139 9132 15476 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15838 9120 15844 9172
rect 15896 9160 15902 9172
rect 16393 9163 16451 9169
rect 16393 9160 16405 9163
rect 15896 9132 16405 9160
rect 15896 9120 15902 9132
rect 16393 9129 16405 9132
rect 16439 9129 16451 9163
rect 16393 9123 16451 9129
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 18046 9160 18052 9172
rect 17635 9132 18052 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 19242 9160 19248 9172
rect 18156 9132 19248 9160
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17092 9064 17816 9092
rect 17092 9052 17098 9064
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 15562 9024 15568 9036
rect 15523 8996 15568 9024
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 9024 15899 9027
rect 15930 9024 15936 9036
rect 15887 8996 15936 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 9024 17187 9027
rect 17494 9024 17500 9036
rect 17175 8996 17500 9024
rect 17175 8993 17187 8996
rect 17129 8987 17187 8993
rect 17494 8984 17500 8996
rect 17552 9024 17558 9036
rect 17788 9024 17816 9064
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 18156 9092 18184 9132
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 20898 9120 20904 9172
rect 20956 9160 20962 9172
rect 21453 9163 21511 9169
rect 21453 9160 21465 9163
rect 20956 9132 21465 9160
rect 20956 9120 20962 9132
rect 21453 9129 21465 9132
rect 21499 9160 21511 9163
rect 21637 9163 21695 9169
rect 21499 9132 21588 9160
rect 21499 9129 21511 9132
rect 21453 9123 21511 9129
rect 18509 9095 18567 9101
rect 18509 9092 18521 9095
rect 17920 9064 18184 9092
rect 18248 9064 18521 9092
rect 17920 9052 17926 9064
rect 18248 9024 18276 9064
rect 18509 9061 18521 9064
rect 18555 9061 18567 9095
rect 18509 9055 18567 9061
rect 19426 9052 19432 9104
rect 19484 9092 19490 9104
rect 19521 9095 19579 9101
rect 19521 9092 19533 9095
rect 19484 9064 19533 9092
rect 19484 9052 19490 9064
rect 19521 9061 19533 9064
rect 19567 9061 19579 9095
rect 19521 9055 19579 9061
rect 17552 8996 17724 9024
rect 17788 8996 18276 9024
rect 18432 8996 21220 9024
rect 17552 8984 17558 8996
rect 3970 8956 3976 8968
rect 3931 8928 3976 8956
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 5810 8956 5816 8968
rect 4663 8928 5816 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 16485 8959 16543 8965
rect 16485 8925 16497 8959
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 1946 8888 1952 8900
rect 1627 8860 1952 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 1946 8848 1952 8860
rect 2004 8848 2010 8900
rect 14826 8848 14832 8900
rect 14884 8848 14890 8900
rect 16500 8888 16528 8919
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17586 8956 17592 8968
rect 17276 8928 17321 8956
rect 17547 8928 17592 8956
rect 17276 8916 17282 8928
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 17696 8956 17724 8996
rect 17954 8956 17960 8968
rect 17696 8928 17960 8956
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18138 8916 18144 8968
rect 18196 8956 18202 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18196 8928 18245 8956
rect 18196 8916 18202 8928
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 16850 8888 16856 8900
rect 16500 8860 16856 8888
rect 16850 8848 16856 8860
rect 16908 8888 16914 8900
rect 17604 8888 17632 8916
rect 17862 8888 17868 8900
rect 16908 8860 17632 8888
rect 17696 8860 17868 8888
rect 16908 8848 16914 8860
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 4338 8820 4344 8832
rect 3927 8792 4344 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 17696 8820 17724 8860
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 18322 8888 18328 8900
rect 18283 8860 18328 8888
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 17184 8792 17724 8820
rect 17773 8823 17831 8829
rect 17184 8780 17190 8792
rect 17773 8789 17785 8823
rect 17819 8820 17831 8823
rect 18432 8820 18460 8996
rect 18782 8916 18788 8968
rect 18840 8956 18846 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 18840 8928 19257 8956
rect 18840 8916 18846 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19978 8916 19984 8968
rect 20036 8956 20042 8968
rect 21192 8965 21220 8996
rect 21266 8984 21272 9036
rect 21324 9024 21330 9036
rect 21560 9024 21588 9132
rect 21637 9129 21649 9163
rect 21683 9160 21695 9163
rect 22094 9160 22100 9172
rect 21683 9132 22100 9160
rect 21683 9129 21695 9132
rect 21637 9123 21695 9129
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22204 9132 22293 9160
rect 22002 9052 22008 9104
rect 22060 9092 22066 9104
rect 22204 9092 22232 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22738 9160 22744 9172
rect 22699 9132 22744 9160
rect 22281 9123 22339 9129
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 23661 9163 23719 9169
rect 23661 9129 23673 9163
rect 23707 9160 23719 9163
rect 25038 9160 25044 9172
rect 23707 9132 25044 9160
rect 23707 9129 23719 9132
rect 23661 9123 23719 9129
rect 25038 9120 25044 9132
rect 25096 9160 25102 9172
rect 29641 9163 29699 9169
rect 29641 9160 29653 9163
rect 25096 9132 29653 9160
rect 25096 9120 25102 9132
rect 29641 9129 29653 9132
rect 29687 9129 29699 9163
rect 29641 9123 29699 9129
rect 30006 9120 30012 9172
rect 30064 9160 30070 9172
rect 31205 9163 31263 9169
rect 31205 9160 31217 9163
rect 30064 9132 31217 9160
rect 30064 9120 30070 9132
rect 31205 9129 31217 9132
rect 31251 9129 31263 9163
rect 35434 9160 35440 9172
rect 35395 9132 35440 9160
rect 31205 9123 31263 9129
rect 35434 9120 35440 9132
rect 35492 9120 35498 9172
rect 22922 9092 22928 9104
rect 22060 9064 22232 9092
rect 22296 9064 22928 9092
rect 22060 9052 22066 9064
rect 22296 9024 22324 9064
rect 22922 9052 22928 9064
rect 22980 9052 22986 9104
rect 23106 9052 23112 9104
rect 23164 9092 23170 9104
rect 24670 9092 24676 9104
rect 23164 9064 24676 9092
rect 23164 9052 23170 9064
rect 24670 9052 24676 9064
rect 24728 9052 24734 9104
rect 24949 9095 25007 9101
rect 24949 9061 24961 9095
rect 24995 9092 25007 9095
rect 25774 9092 25780 9104
rect 24995 9064 25780 9092
rect 24995 9061 25007 9064
rect 24949 9055 25007 9061
rect 25774 9052 25780 9064
rect 25832 9092 25838 9104
rect 26050 9092 26056 9104
rect 25832 9064 26056 9092
rect 25832 9052 25838 9064
rect 26050 9052 26056 9064
rect 26108 9052 26114 9104
rect 27430 9052 27436 9104
rect 27488 9092 27494 9104
rect 27488 9064 28120 9092
rect 27488 9052 27494 9064
rect 24486 9024 24492 9036
rect 21324 8996 21369 9024
rect 21560 8996 22324 9024
rect 22480 8996 24492 9024
rect 21324 8984 21330 8996
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 20036 8928 20177 8956
rect 20036 8916 20042 8928
rect 20165 8925 20177 8928
rect 20211 8925 20223 8959
rect 20165 8919 20223 8925
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8925 21235 8959
rect 21450 8956 21456 8968
rect 21411 8928 21456 8956
rect 21177 8919 21235 8925
rect 21450 8916 21456 8928
rect 21508 8956 21514 8968
rect 22186 8956 22192 8968
rect 21508 8928 22094 8956
rect 22147 8928 22192 8956
rect 21508 8916 21514 8928
rect 18509 8891 18567 8897
rect 18509 8857 18521 8891
rect 18555 8888 18567 8891
rect 19521 8891 19579 8897
rect 18555 8860 19472 8888
rect 18555 8857 18567 8860
rect 18509 8851 18567 8857
rect 17819 8792 18460 8820
rect 17819 8789 17831 8792
rect 17773 8783 17831 8789
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 19337 8823 19395 8829
rect 19337 8820 19349 8823
rect 18932 8792 19349 8820
rect 18932 8780 18938 8792
rect 19337 8789 19349 8792
rect 19383 8789 19395 8823
rect 19444 8820 19472 8860
rect 19521 8857 19533 8891
rect 19567 8888 19579 8891
rect 20622 8888 20628 8900
rect 19567 8860 20628 8888
rect 19567 8857 19579 8860
rect 19521 8851 19579 8857
rect 20622 8848 20628 8860
rect 20680 8848 20686 8900
rect 22066 8888 22094 8928
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 22278 8916 22284 8968
rect 22336 8956 22342 8968
rect 22480 8956 22508 8996
rect 22336 8928 22508 8956
rect 22557 8959 22615 8965
rect 22336 8916 22342 8928
rect 22557 8925 22569 8959
rect 22603 8956 22615 8959
rect 22830 8956 22836 8968
rect 22603 8928 22836 8956
rect 22603 8925 22615 8928
rect 22557 8919 22615 8925
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 23676 8965 23704 8996
rect 24486 8984 24492 8996
rect 24544 8984 24550 9036
rect 25038 9024 25044 9036
rect 24596 8996 25044 9024
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24596 8956 24624 8996
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 25590 8984 25596 9036
rect 25648 9024 25654 9036
rect 25961 9027 26019 9033
rect 25961 9024 25973 9027
rect 25648 8996 25973 9024
rect 25648 8984 25654 8996
rect 25961 8993 25973 8996
rect 26007 8993 26019 9027
rect 25961 8987 26019 8993
rect 26245 9027 26303 9033
rect 26245 8993 26257 9027
rect 26291 9024 26303 9027
rect 26418 9024 26424 9036
rect 26291 8996 26424 9024
rect 26291 8993 26303 8996
rect 26245 8987 26303 8993
rect 26418 8984 26424 8996
rect 26476 8984 26482 9036
rect 28092 9024 28120 9064
rect 28534 9052 28540 9104
rect 28592 9092 28598 9104
rect 30561 9095 30619 9101
rect 30561 9092 30573 9095
rect 28592 9064 30573 9092
rect 28592 9052 28598 9064
rect 30561 9061 30573 9064
rect 30607 9061 30619 9095
rect 30561 9055 30619 9061
rect 37182 9024 37188 9036
rect 28092 8996 29592 9024
rect 37143 8996 37188 9024
rect 25130 8956 25136 8968
rect 23891 8928 24624 8956
rect 24688 8928 25136 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 22462 8888 22468 8900
rect 21560 8860 21772 8888
rect 22066 8860 22468 8888
rect 20070 8820 20076 8832
rect 19444 8792 20076 8820
rect 19337 8783 19395 8789
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 20257 8823 20315 8829
rect 20257 8789 20269 8823
rect 20303 8820 20315 8823
rect 21560 8820 21588 8860
rect 20303 8792 21588 8820
rect 21744 8820 21772 8860
rect 22462 8848 22468 8860
rect 22520 8848 22526 8900
rect 24581 8891 24639 8897
rect 24581 8857 24593 8891
rect 24627 8888 24639 8891
rect 24688 8888 24716 8928
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 26050 8956 26056 8968
rect 26011 8928 26056 8956
rect 26050 8916 26056 8928
rect 26108 8916 26114 8968
rect 26145 8959 26203 8965
rect 26145 8925 26157 8959
rect 26191 8925 26203 8959
rect 26145 8919 26203 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 27798 8956 27804 8968
rect 27203 8928 27804 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 24627 8860 24716 8888
rect 24627 8857 24639 8860
rect 24581 8851 24639 8857
rect 24762 8848 24768 8900
rect 24820 8888 24826 8900
rect 24820 8860 24865 8888
rect 24820 8848 24826 8860
rect 22738 8820 22744 8832
rect 21744 8792 22744 8820
rect 20303 8789 20315 8792
rect 20257 8783 20315 8789
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 24394 8820 24400 8832
rect 24355 8792 24400 8820
rect 24394 8780 24400 8792
rect 24452 8780 24458 8832
rect 24670 8780 24676 8832
rect 24728 8820 24734 8832
rect 26160 8820 26188 8919
rect 27798 8916 27804 8928
rect 27856 8956 27862 8968
rect 27893 8959 27951 8965
rect 27893 8956 27905 8959
rect 27856 8928 27905 8956
rect 27856 8916 27862 8928
rect 27893 8925 27905 8928
rect 27939 8925 27951 8959
rect 27893 8919 27951 8925
rect 28169 8959 28227 8965
rect 28169 8925 28181 8959
rect 28215 8956 28227 8959
rect 28258 8956 28264 8968
rect 28215 8928 28264 8956
rect 28215 8925 28227 8928
rect 28169 8919 28227 8925
rect 28258 8916 28264 8928
rect 28316 8916 28322 8968
rect 29564 8965 29592 8996
rect 37182 8984 37188 8996
rect 37240 8984 37246 9036
rect 37918 9024 37924 9036
rect 37879 8996 37924 9024
rect 37918 8984 37924 8996
rect 37976 8984 37982 9036
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 29638 8916 29644 8968
rect 29696 8956 29702 8968
rect 29825 8959 29883 8965
rect 29825 8956 29837 8959
rect 29696 8928 29837 8956
rect 29696 8916 29702 8928
rect 29825 8925 29837 8928
rect 29871 8956 29883 8959
rect 30190 8956 30196 8968
rect 29871 8928 30196 8956
rect 29871 8925 29883 8928
rect 29825 8919 29883 8925
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 30374 8916 30380 8968
rect 30432 8956 30438 8968
rect 30653 8959 30711 8965
rect 30653 8956 30665 8959
rect 30432 8928 30665 8956
rect 30432 8916 30438 8928
rect 30653 8925 30665 8928
rect 30699 8956 30711 8959
rect 31113 8959 31171 8965
rect 31113 8956 31125 8959
rect 30699 8928 31125 8956
rect 30699 8925 30711 8928
rect 30653 8919 30711 8925
rect 31113 8925 31125 8928
rect 31159 8925 31171 8959
rect 31113 8919 31171 8925
rect 38102 8916 38108 8968
rect 38160 8956 38166 8968
rect 38160 8928 38205 8956
rect 38160 8916 38166 8928
rect 26878 8888 26884 8900
rect 26839 8860 26884 8888
rect 26878 8848 26884 8860
rect 26936 8848 26942 8900
rect 27065 8891 27123 8897
rect 27065 8857 27077 8891
rect 27111 8888 27123 8891
rect 27111 8860 27384 8888
rect 27111 8857 27123 8860
rect 27065 8851 27123 8857
rect 26234 8820 26240 8832
rect 24728 8792 24773 8820
rect 26160 8792 26240 8820
rect 24728 8780 24734 8792
rect 26234 8780 26240 8792
rect 26292 8780 26298 8832
rect 26418 8820 26424 8832
rect 26379 8792 26424 8820
rect 26418 8780 26424 8792
rect 26476 8780 26482 8832
rect 26786 8780 26792 8832
rect 26844 8820 26850 8832
rect 27249 8823 27307 8829
rect 27249 8820 27261 8823
rect 26844 8792 27261 8820
rect 26844 8780 26850 8792
rect 27249 8789 27261 8792
rect 27295 8789 27307 8823
rect 27356 8820 27384 8860
rect 27430 8848 27436 8900
rect 27488 8888 27494 8900
rect 27488 8860 27533 8888
rect 27488 8848 27494 8860
rect 27982 8848 27988 8900
rect 28040 8888 28046 8900
rect 30009 8891 30067 8897
rect 30009 8888 30021 8891
rect 28040 8860 30021 8888
rect 28040 8848 28046 8860
rect 30009 8857 30021 8860
rect 30055 8857 30067 8891
rect 30009 8851 30067 8857
rect 27614 8820 27620 8832
rect 27356 8792 27620 8820
rect 27249 8783 27307 8789
rect 27614 8780 27620 8792
rect 27672 8820 27678 8832
rect 28074 8820 28080 8832
rect 27672 8792 28080 8820
rect 27672 8780 27678 8792
rect 28074 8780 28080 8792
rect 28132 8780 28138 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 13596 8588 14841 8616
rect 13596 8576 13602 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 16666 8616 16672 8628
rect 16627 8588 16672 8616
rect 14829 8579 14887 8585
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 17460 8588 17969 8616
rect 17460 8576 17466 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18230 8616 18236 8628
rect 18187 8588 18236 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 20404 8588 20453 8616
rect 20404 8576 20410 8588
rect 20441 8585 20453 8588
rect 20487 8616 20499 8619
rect 22830 8616 22836 8628
rect 20487 8588 21128 8616
rect 22791 8588 22836 8616
rect 20487 8585 20499 8588
rect 20441 8579 20499 8585
rect 4338 8548 4344 8560
rect 4299 8520 4344 8548
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 18782 8557 18788 8560
rect 17773 8551 17831 8557
rect 17773 8548 17785 8551
rect 17696 8520 17785 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2130 8480 2136 8492
rect 2087 8452 2136 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 7926 8480 7932 8492
rect 5215 8452 7932 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 7926 8440 7932 8452
rect 7984 8480 7990 8492
rect 9950 8480 9956 8492
rect 7984 8452 9956 8480
rect 7984 8440 7990 8452
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 15194 8480 15200 8492
rect 15155 8452 15200 8480
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 16850 8480 16856 8492
rect 16811 8452 16856 8480
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 17184 8452 17229 8480
rect 17184 8440 17190 8452
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 17696 8480 17724 8520
rect 17773 8517 17785 8520
rect 17819 8517 17831 8551
rect 17773 8511 17831 8517
rect 18769 8551 18788 8557
rect 18769 8517 18781 8551
rect 18769 8511 18788 8517
rect 18782 8508 18788 8511
rect 18840 8508 18846 8560
rect 18969 8551 19027 8557
rect 18969 8517 18981 8551
rect 19015 8548 19027 8551
rect 19058 8548 19064 8560
rect 19015 8520 19064 8548
rect 19015 8517 19027 8520
rect 18969 8511 19027 8517
rect 19058 8508 19064 8520
rect 19116 8508 19122 8560
rect 19426 8508 19432 8560
rect 19484 8548 19490 8560
rect 21100 8557 21128 8588
rect 22830 8576 22836 8588
rect 22888 8576 22894 8628
rect 23934 8616 23940 8628
rect 23895 8588 23940 8616
rect 23934 8576 23940 8588
rect 23992 8576 23998 8628
rect 24305 8619 24363 8625
rect 24305 8585 24317 8619
rect 24351 8616 24363 8619
rect 24670 8616 24676 8628
rect 24351 8588 24676 8616
rect 24351 8585 24363 8588
rect 24305 8579 24363 8585
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 24854 8616 24860 8628
rect 24815 8588 24860 8616
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 26878 8616 26884 8628
rect 25188 8588 26884 8616
rect 25188 8576 25194 8588
rect 26878 8576 26884 8588
rect 26936 8576 26942 8628
rect 27798 8576 27804 8628
rect 27856 8616 27862 8628
rect 29638 8616 29644 8628
rect 27856 8588 29644 8616
rect 27856 8576 27862 8588
rect 29638 8576 29644 8588
rect 29696 8576 29702 8628
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 19484 8520 19809 8548
rect 19484 8508 19490 8520
rect 19797 8517 19809 8520
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 21085 8551 21143 8557
rect 21085 8517 21097 8551
rect 21131 8517 21143 8551
rect 23106 8548 23112 8560
rect 21085 8511 21143 8517
rect 21284 8520 23112 8548
rect 17552 8452 17724 8480
rect 17552 8440 17558 8452
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 17920 8452 17965 8480
rect 17920 8440 17926 8452
rect 19334 8440 19340 8492
rect 19392 8480 19398 8492
rect 19613 8483 19671 8489
rect 19392 8452 19564 8480
rect 19392 8440 19398 8452
rect 2866 8412 2872 8424
rect 2827 8384 2872 8412
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 4120 8384 4537 8412
rect 4120 8372 4126 8384
rect 4525 8381 4537 8384
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 15289 8415 15347 8421
rect 15289 8381 15301 8415
rect 15335 8412 15347 8415
rect 15378 8412 15384 8424
rect 15335 8384 15384 8412
rect 15335 8381 15347 8384
rect 15289 8375 15347 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15654 8412 15660 8424
rect 15519 8384 15660 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15654 8372 15660 8384
rect 15712 8412 15718 8424
rect 19429 8415 19487 8421
rect 19429 8412 19441 8415
rect 15712 8384 16896 8412
rect 15712 8372 15718 8384
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5626 8344 5632 8356
rect 5123 8316 5632 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 16868 8276 16896 8384
rect 17236 8384 19441 8412
rect 16942 8304 16948 8356
rect 17000 8344 17006 8356
rect 17236 8344 17264 8384
rect 19429 8381 19441 8384
rect 19475 8381 19487 8415
rect 19536 8412 19564 8452
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 20070 8480 20076 8492
rect 19659 8452 20076 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 20070 8440 20076 8452
rect 20128 8480 20134 8492
rect 20349 8483 20407 8489
rect 20349 8480 20361 8483
rect 20128 8452 20361 8480
rect 20128 8440 20134 8452
rect 20349 8449 20361 8452
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 20530 8440 20536 8492
rect 20588 8480 20594 8492
rect 21174 8480 21180 8492
rect 20588 8452 21180 8480
rect 20588 8440 20594 8452
rect 21174 8440 21180 8452
rect 21232 8480 21238 8492
rect 21284 8489 21312 8520
rect 23106 8508 23112 8520
rect 23164 8508 23170 8560
rect 23198 8508 23204 8560
rect 23256 8548 23262 8560
rect 23753 8551 23811 8557
rect 23753 8548 23765 8551
rect 23256 8520 23765 8548
rect 23256 8508 23262 8520
rect 23753 8517 23765 8520
rect 23799 8517 23811 8551
rect 23753 8511 23811 8517
rect 24029 8551 24087 8557
rect 24029 8517 24041 8551
rect 24075 8548 24087 8551
rect 25038 8548 25044 8560
rect 24075 8520 24808 8548
rect 24951 8520 25044 8548
rect 24075 8517 24087 8520
rect 24029 8511 24087 8517
rect 24780 8492 24808 8520
rect 25038 8508 25044 8520
rect 25096 8548 25102 8560
rect 25096 8520 26188 8548
rect 25096 8508 25102 8520
rect 21269 8483 21327 8489
rect 21269 8480 21281 8483
rect 21232 8452 21281 8480
rect 21232 8440 21238 8452
rect 21269 8449 21281 8452
rect 21315 8449 21327 8483
rect 22002 8480 22008 8492
rect 21963 8452 22008 8480
rect 21269 8443 21327 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 22741 8483 22799 8489
rect 22741 8449 22753 8483
rect 22787 8480 22799 8483
rect 22830 8480 22836 8492
rect 22787 8452 22836 8480
rect 22787 8449 22799 8452
rect 22741 8443 22799 8449
rect 22830 8440 22836 8452
rect 22888 8440 22894 8492
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8480 22983 8483
rect 23290 8480 23296 8492
rect 22971 8452 23296 8480
rect 22971 8449 22983 8452
rect 22925 8443 22983 8449
rect 23290 8440 23296 8452
rect 23348 8440 23354 8492
rect 24121 8483 24179 8489
rect 24121 8449 24133 8483
rect 24167 8449 24179 8483
rect 24762 8480 24768 8492
rect 24723 8452 24768 8480
rect 24121 8443 24179 8449
rect 23842 8412 23848 8424
rect 19536 8384 23848 8412
rect 19429 8375 19487 8381
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 24136 8412 24164 8443
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 25130 8480 25136 8492
rect 25091 8452 25136 8480
rect 25130 8440 25136 8452
rect 25188 8440 25194 8492
rect 26160 8489 26188 8520
rect 26418 8508 26424 8560
rect 26476 8548 26482 8560
rect 28997 8551 29055 8557
rect 28997 8548 29009 8551
rect 26476 8520 29009 8548
rect 26476 8508 26482 8520
rect 28997 8517 29009 8520
rect 29043 8517 29055 8551
rect 30926 8548 30932 8560
rect 30222 8520 30932 8548
rect 28997 8511 29055 8517
rect 30926 8508 30932 8520
rect 30984 8508 30990 8560
rect 26145 8483 26203 8489
rect 26145 8449 26157 8483
rect 26191 8480 26203 8483
rect 26326 8480 26332 8492
rect 26191 8452 26332 8480
rect 26191 8449 26203 8452
rect 26145 8443 26203 8449
rect 26326 8440 26332 8452
rect 26384 8440 26390 8492
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8480 27491 8483
rect 27614 8480 27620 8492
rect 27479 8452 27620 8480
rect 27479 8449 27491 8452
rect 27433 8443 27491 8449
rect 27614 8440 27620 8452
rect 27672 8440 27678 8492
rect 36722 8480 36728 8492
rect 36683 8452 36728 8480
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 37829 8483 37887 8489
rect 37829 8449 37841 8483
rect 37875 8480 37887 8483
rect 38102 8480 38108 8492
rect 37875 8452 38108 8480
rect 37875 8449 37887 8452
rect 37829 8443 37887 8449
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 24949 8415 25007 8421
rect 24949 8412 24961 8415
rect 24136 8384 24961 8412
rect 24949 8381 24961 8384
rect 24995 8412 25007 8415
rect 25222 8412 25228 8424
rect 24995 8384 25228 8412
rect 24995 8381 25007 8384
rect 24949 8375 25007 8381
rect 25222 8372 25228 8384
rect 25280 8372 25286 8424
rect 26418 8412 26424 8424
rect 26379 8384 26424 8412
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 27709 8415 27767 8421
rect 27709 8412 27721 8415
rect 27264 8384 27721 8412
rect 17000 8316 17264 8344
rect 17589 8347 17647 8353
rect 17000 8304 17006 8316
rect 17589 8313 17601 8347
rect 17635 8344 17647 8347
rect 18046 8344 18052 8356
rect 17635 8316 18052 8344
rect 17635 8313 17647 8316
rect 17589 8307 17647 8313
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 18230 8304 18236 8356
rect 18288 8344 18294 8356
rect 18288 8316 18828 8344
rect 18288 8304 18294 8316
rect 18800 8285 18828 8316
rect 20622 8304 20628 8356
rect 20680 8344 20686 8356
rect 23750 8344 23756 8356
rect 20680 8316 23756 8344
rect 20680 8304 20686 8316
rect 23750 8304 23756 8316
rect 23808 8344 23814 8356
rect 24302 8344 24308 8356
rect 23808 8316 24308 8344
rect 23808 8304 23814 8316
rect 24302 8304 24308 8316
rect 24360 8304 24366 8356
rect 25866 8304 25872 8356
rect 25924 8344 25930 8356
rect 27264 8344 27292 8384
rect 27709 8381 27721 8384
rect 27755 8412 27767 8415
rect 27798 8412 27804 8424
rect 27755 8384 27804 8412
rect 27755 8381 27767 8384
rect 27709 8375 27767 8381
rect 27798 8372 27804 8384
rect 27856 8372 27862 8424
rect 28718 8412 28724 8424
rect 28679 8384 28724 8412
rect 28718 8372 28724 8384
rect 28776 8372 28782 8424
rect 30469 8415 30527 8421
rect 30469 8412 30481 8415
rect 28828 8384 30481 8412
rect 25924 8316 27292 8344
rect 25924 8304 25930 8316
rect 27614 8304 27620 8356
rect 27672 8344 27678 8356
rect 28828 8344 28856 8384
rect 30469 8381 30481 8384
rect 30515 8381 30527 8415
rect 30469 8375 30527 8381
rect 27672 8316 28856 8344
rect 27672 8304 27678 8316
rect 18601 8279 18659 8285
rect 18601 8276 18613 8279
rect 16868 8248 18613 8276
rect 18601 8245 18613 8248
rect 18647 8245 18659 8279
rect 18601 8239 18659 8245
rect 18785 8279 18843 8285
rect 18785 8245 18797 8279
rect 18831 8245 18843 8279
rect 18785 8239 18843 8245
rect 22189 8279 22247 8285
rect 22189 8245 22201 8279
rect 22235 8276 22247 8279
rect 22370 8276 22376 8288
rect 22235 8248 22376 8276
rect 22235 8245 22247 8248
rect 22189 8239 22247 8245
rect 22370 8236 22376 8248
rect 22428 8236 22434 8288
rect 23474 8236 23480 8288
rect 23532 8276 23538 8288
rect 24026 8276 24032 8288
rect 23532 8248 24032 8276
rect 23532 8236 23538 8248
rect 24026 8236 24032 8248
rect 24084 8236 24090 8288
rect 24762 8236 24768 8288
rect 24820 8276 24826 8288
rect 25314 8276 25320 8288
rect 24820 8248 25320 8276
rect 24820 8236 24826 8248
rect 25314 8236 25320 8248
rect 25372 8236 25378 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 15252 8044 15485 8072
rect 15252 8032 15258 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 15473 8035 15531 8041
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18417 8075 18475 8081
rect 18417 8072 18429 8075
rect 18196 8044 18429 8072
rect 18196 8032 18202 8044
rect 18417 8041 18429 8044
rect 18463 8041 18475 8075
rect 18417 8035 18475 8041
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 18564 8044 19625 8072
rect 18564 8032 18570 8044
rect 19613 8041 19625 8044
rect 19659 8072 19671 8075
rect 22189 8075 22247 8081
rect 19659 8044 21680 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 2130 7964 2136 8016
rect 2188 8004 2194 8016
rect 17405 8007 17463 8013
rect 2188 7976 6914 8004
rect 2188 7964 2194 7976
rect 3970 7936 3976 7948
rect 3931 7908 3976 7936
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 5626 7936 5632 7948
rect 5587 7908 5632 7936
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6886 7936 6914 7976
rect 17405 7973 17417 8007
rect 17451 8004 17463 8007
rect 18782 8004 18788 8016
rect 17451 7976 18788 8004
rect 17451 7973 17463 7976
rect 17405 7967 17463 7973
rect 18782 7964 18788 7976
rect 18840 7964 18846 8016
rect 21450 8004 21456 8016
rect 18892 7976 21456 8004
rect 18892 7936 18920 7976
rect 21450 7964 21456 7976
rect 21508 7964 21514 8016
rect 6886 7908 18920 7936
rect 21652 7936 21680 8044
rect 22189 8041 22201 8075
rect 22235 8072 22247 8075
rect 22646 8072 22652 8084
rect 22235 8044 22652 8072
rect 22235 8041 22247 8044
rect 22189 8035 22247 8041
rect 22646 8032 22652 8044
rect 22704 8032 22710 8084
rect 23661 8075 23719 8081
rect 23661 8041 23673 8075
rect 23707 8072 23719 8075
rect 25038 8072 25044 8084
rect 23707 8044 25044 8072
rect 23707 8041 23719 8044
rect 23661 8035 23719 8041
rect 25038 8032 25044 8044
rect 25096 8032 25102 8084
rect 26050 8032 26056 8084
rect 26108 8072 26114 8084
rect 30285 8075 30343 8081
rect 30285 8072 30297 8075
rect 26108 8044 30297 8072
rect 26108 8032 26114 8044
rect 30285 8041 30297 8044
rect 30331 8041 30343 8075
rect 30926 8072 30932 8084
rect 30887 8044 30932 8072
rect 30285 8035 30343 8041
rect 30926 8032 30932 8044
rect 30984 8032 30990 8084
rect 38010 8032 38016 8084
rect 38068 8072 38074 8084
rect 38105 8075 38163 8081
rect 38105 8072 38117 8075
rect 38068 8044 38117 8072
rect 38068 8032 38074 8044
rect 38105 8041 38117 8044
rect 38151 8041 38163 8075
rect 38105 8035 38163 8041
rect 22094 7964 22100 8016
rect 22152 8004 22158 8016
rect 22925 8007 22983 8013
rect 22925 8004 22937 8007
rect 22152 7976 22937 8004
rect 22152 7964 22158 7976
rect 22925 7973 22937 7976
rect 22971 7973 22983 8007
rect 22925 7967 22983 7973
rect 23845 8007 23903 8013
rect 23845 7973 23857 8007
rect 23891 8004 23903 8007
rect 25498 8004 25504 8016
rect 23891 7976 25504 8004
rect 23891 7973 23903 7976
rect 23845 7967 23903 7973
rect 25498 7964 25504 7976
rect 25556 7964 25562 8016
rect 25866 7964 25872 8016
rect 25924 8004 25930 8016
rect 25924 7976 26188 8004
rect 25924 7964 25930 7976
rect 22186 7936 22192 7948
rect 21652 7908 22192 7936
rect 22186 7896 22192 7908
rect 22244 7896 22250 7948
rect 26160 7945 26188 7976
rect 26418 7964 26424 8016
rect 26476 8004 26482 8016
rect 27522 8004 27528 8016
rect 26476 7976 27528 8004
rect 26476 7964 26482 7976
rect 27522 7964 27528 7976
rect 27580 7964 27586 8016
rect 27798 7964 27804 8016
rect 27856 8004 27862 8016
rect 27856 7976 35020 8004
rect 27856 7964 27862 7976
rect 26145 7939 26203 7945
rect 26145 7905 26157 7939
rect 26191 7905 26203 7939
rect 26145 7899 26203 7905
rect 26237 7939 26295 7945
rect 26237 7905 26249 7939
rect 26283 7936 26295 7939
rect 26326 7936 26332 7948
rect 26283 7908 26332 7936
rect 26283 7905 26295 7908
rect 26237 7899 26295 7905
rect 26326 7896 26332 7908
rect 26384 7896 26390 7948
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 15378 7868 15384 7880
rect 15339 7840 15384 7868
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7868 15623 7871
rect 15746 7868 15752 7880
rect 15611 7840 15752 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7837 16267 7871
rect 16390 7868 16396 7880
rect 16351 7840 16396 7868
rect 16209 7831 16267 7837
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 16025 7735 16083 7741
rect 16025 7732 16037 7735
rect 15804 7704 16037 7732
rect 15804 7692 15810 7704
rect 16025 7701 16037 7704
rect 16071 7701 16083 7735
rect 16224 7732 16252 7831
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 17034 7868 17040 7880
rect 16995 7840 17040 7868
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 17267 7840 18245 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 18233 7837 18245 7840
rect 18279 7868 18291 7871
rect 18690 7868 18696 7880
rect 18279 7840 18696 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18690 7828 18696 7840
rect 18748 7868 18754 7880
rect 20806 7868 20812 7880
rect 18748 7840 19564 7868
rect 18748 7828 18754 7840
rect 17862 7800 17868 7812
rect 17823 7772 17868 7800
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 17954 7760 17960 7812
rect 18012 7800 18018 7812
rect 18049 7803 18107 7809
rect 18049 7800 18061 7803
rect 18012 7772 18061 7800
rect 18012 7760 18018 7772
rect 18049 7769 18061 7772
rect 18095 7769 18107 7803
rect 18049 7763 18107 7769
rect 18141 7803 18199 7809
rect 18141 7769 18153 7803
rect 18187 7800 18199 7803
rect 19334 7800 19340 7812
rect 18187 7772 19340 7800
rect 18187 7769 18199 7772
rect 18141 7763 18199 7769
rect 19334 7760 19340 7772
rect 19392 7760 19398 7812
rect 18230 7732 18236 7744
rect 16224 7704 18236 7732
rect 16025 7695 16083 7701
rect 18230 7692 18236 7704
rect 18288 7732 18294 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 18288 7704 19441 7732
rect 18288 7692 18294 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 19536 7732 19564 7840
rect 19720 7840 20812 7868
rect 19597 7803 19655 7809
rect 19597 7769 19609 7803
rect 19643 7800 19655 7803
rect 19720 7800 19748 7840
rect 20806 7828 20812 7840
rect 20864 7868 20870 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20864 7840 20913 7868
rect 20864 7828 20870 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7837 21235 7871
rect 22370 7868 22376 7880
rect 22331 7840 22376 7868
rect 21177 7831 21235 7837
rect 19643 7772 19748 7800
rect 19797 7803 19855 7809
rect 19643 7769 19655 7772
rect 19597 7763 19655 7769
rect 19797 7769 19809 7803
rect 19843 7800 19855 7803
rect 20714 7800 20720 7812
rect 19843 7772 20720 7800
rect 19843 7769 19855 7772
rect 19797 7763 19855 7769
rect 20714 7760 20720 7772
rect 20772 7800 20778 7812
rect 20990 7800 20996 7812
rect 20772 7772 20996 7800
rect 20772 7760 20778 7772
rect 20990 7760 20996 7772
rect 21048 7760 21054 7812
rect 21192 7800 21220 7831
rect 22370 7828 22376 7840
rect 22428 7828 22434 7880
rect 24394 7868 24400 7880
rect 22848 7840 24400 7868
rect 22848 7800 22876 7840
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7868 25007 7871
rect 25130 7868 25136 7880
rect 24995 7840 25136 7868
rect 24995 7837 25007 7840
rect 24949 7831 25007 7837
rect 21192 7772 22876 7800
rect 21192 7732 21220 7772
rect 22922 7760 22928 7812
rect 22980 7800 22986 7812
rect 23382 7800 23388 7812
rect 22980 7772 23388 7800
rect 22980 7760 22986 7772
rect 23382 7760 23388 7772
rect 23440 7760 23446 7812
rect 23474 7760 23480 7812
rect 23532 7800 23538 7812
rect 23693 7803 23751 7809
rect 23532 7772 23577 7800
rect 23532 7760 23538 7772
rect 23693 7769 23705 7803
rect 23739 7800 23751 7803
rect 24964 7800 24992 7831
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 25682 7828 25688 7880
rect 25740 7868 25746 7880
rect 25961 7871 26019 7877
rect 25961 7868 25973 7871
rect 25740 7840 25973 7868
rect 25740 7828 25746 7840
rect 25961 7837 25973 7840
rect 26007 7837 26019 7871
rect 25961 7831 26019 7837
rect 23739 7772 24992 7800
rect 23739 7769 23751 7772
rect 23693 7763 23751 7769
rect 25038 7760 25044 7812
rect 25096 7800 25102 7812
rect 25314 7800 25320 7812
rect 25096 7772 25141 7800
rect 25275 7772 25320 7800
rect 25096 7760 25102 7772
rect 25314 7760 25320 7772
rect 25372 7760 25378 7812
rect 19536 7704 21220 7732
rect 22465 7735 22523 7741
rect 19429 7695 19487 7701
rect 22465 7701 22477 7735
rect 22511 7732 22523 7735
rect 23842 7732 23848 7744
rect 22511 7704 23848 7732
rect 22511 7701 22523 7704
rect 22465 7695 22523 7701
rect 23842 7692 23848 7704
rect 23900 7692 23906 7744
rect 24762 7732 24768 7744
rect 24723 7704 24768 7732
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 25133 7735 25191 7741
rect 25133 7701 25145 7735
rect 25179 7732 25191 7735
rect 25222 7732 25228 7744
rect 25179 7704 25228 7732
rect 25179 7701 25191 7704
rect 25133 7695 25191 7701
rect 25222 7692 25228 7704
rect 25280 7692 25286 7744
rect 25976 7732 26004 7831
rect 26050 7828 26056 7880
rect 26108 7868 26114 7880
rect 26881 7871 26939 7877
rect 26108 7840 26153 7868
rect 26108 7828 26114 7840
rect 26881 7837 26893 7871
rect 26927 7837 26939 7871
rect 26881 7831 26939 7837
rect 26786 7800 26792 7812
rect 26344 7772 26792 7800
rect 26344 7732 26372 7772
rect 26786 7760 26792 7772
rect 26844 7800 26850 7812
rect 26896 7800 26924 7831
rect 26970 7828 26976 7880
rect 27028 7877 27034 7880
rect 27028 7871 27077 7877
rect 27028 7837 27031 7871
rect 27065 7837 27077 7871
rect 27028 7831 27077 7837
rect 27028 7828 27034 7831
rect 27154 7828 27160 7880
rect 27212 7868 27218 7880
rect 27341 7871 27399 7877
rect 27212 7840 27257 7868
rect 27212 7828 27218 7840
rect 27341 7837 27353 7871
rect 27387 7868 27399 7871
rect 27387 7840 27476 7868
rect 27387 7837 27399 7840
rect 27341 7831 27399 7837
rect 27246 7800 27252 7812
rect 26844 7772 26924 7800
rect 27207 7772 27252 7800
rect 26844 7760 26850 7772
rect 27246 7760 27252 7772
rect 27304 7760 27310 7812
rect 25976 7704 26372 7732
rect 26421 7735 26479 7741
rect 26421 7701 26433 7735
rect 26467 7732 26479 7735
rect 27448 7732 27476 7840
rect 27522 7828 27528 7880
rect 27580 7868 27586 7880
rect 28169 7871 28227 7877
rect 27580 7840 28120 7868
rect 27580 7828 27586 7840
rect 27798 7800 27804 7812
rect 27540 7772 27804 7800
rect 27540 7741 27568 7772
rect 27798 7760 27804 7772
rect 27856 7760 27862 7812
rect 27890 7760 27896 7812
rect 27948 7800 27954 7812
rect 27985 7803 28043 7809
rect 27985 7800 27997 7803
rect 27948 7772 27997 7800
rect 27948 7760 27954 7772
rect 27985 7769 27997 7772
rect 28031 7769 28043 7803
rect 28092 7800 28120 7840
rect 28169 7837 28181 7871
rect 28215 7868 28227 7871
rect 28258 7868 28264 7880
rect 28215 7840 28264 7868
rect 28215 7837 28227 7840
rect 28169 7831 28227 7837
rect 28258 7828 28264 7840
rect 28316 7828 28322 7880
rect 28353 7871 28411 7877
rect 28353 7837 28365 7871
rect 28399 7837 28411 7871
rect 28353 7831 28411 7837
rect 28537 7871 28595 7877
rect 28537 7837 28549 7871
rect 28583 7868 28595 7871
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 28583 7840 29561 7868
rect 28583 7837 28595 7840
rect 28537 7831 28595 7837
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 30190 7868 30196 7880
rect 30151 7840 30196 7868
rect 29549 7831 29607 7837
rect 28368 7800 28396 7831
rect 30190 7828 30196 7840
rect 30248 7828 30254 7880
rect 30374 7828 30380 7880
rect 30432 7868 30438 7880
rect 34992 7877 35020 7976
rect 31021 7871 31079 7877
rect 31021 7868 31033 7871
rect 30432 7840 31033 7868
rect 30432 7828 30438 7840
rect 31021 7837 31033 7840
rect 31067 7837 31079 7871
rect 31021 7831 31079 7837
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7837 35035 7871
rect 35618 7868 35624 7880
rect 35579 7840 35624 7868
rect 34977 7831 35035 7837
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 28092 7772 28396 7800
rect 27985 7763 28043 7769
rect 28442 7760 28448 7812
rect 28500 7800 28506 7812
rect 29641 7803 29699 7809
rect 29641 7800 29653 7803
rect 28500 7772 29653 7800
rect 28500 7760 28506 7772
rect 29641 7769 29653 7772
rect 29687 7769 29699 7803
rect 29641 7763 29699 7769
rect 35069 7803 35127 7809
rect 35069 7769 35081 7803
rect 35115 7800 35127 7803
rect 35805 7803 35863 7809
rect 35805 7800 35817 7803
rect 35115 7772 35817 7800
rect 35115 7769 35127 7772
rect 35069 7763 35127 7769
rect 35805 7769 35817 7772
rect 35851 7769 35863 7803
rect 35805 7763 35863 7769
rect 37461 7803 37519 7809
rect 37461 7769 37473 7803
rect 37507 7800 37519 7803
rect 38654 7800 38660 7812
rect 37507 7772 38660 7800
rect 37507 7769 37519 7772
rect 37461 7763 37519 7769
rect 38654 7760 38660 7772
rect 38712 7760 38718 7812
rect 26467 7704 27476 7732
rect 27525 7735 27583 7741
rect 26467 7701 26479 7704
rect 26421 7695 26479 7701
rect 27525 7701 27537 7735
rect 27571 7701 27583 7735
rect 27525 7695 27583 7701
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 28261 7735 28319 7741
rect 28261 7732 28273 7735
rect 27672 7704 28273 7732
rect 27672 7692 27678 7704
rect 28261 7701 28273 7704
rect 28307 7701 28319 7735
rect 28261 7695 28319 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 15746 7528 15752 7540
rect 15707 7500 15752 7528
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16390 7488 16396 7540
rect 16448 7528 16454 7540
rect 18414 7528 18420 7540
rect 16448 7500 18420 7528
rect 16448 7488 16454 7500
rect 18414 7488 18420 7500
rect 18472 7528 18478 7540
rect 18874 7528 18880 7540
rect 18472 7500 18880 7528
rect 18472 7488 18478 7500
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 20070 7528 20076 7540
rect 20031 7500 20076 7528
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 22186 7528 22192 7540
rect 22147 7500 22192 7528
rect 22186 7488 22192 7500
rect 22244 7488 22250 7540
rect 23385 7531 23443 7537
rect 23385 7497 23397 7531
rect 23431 7528 23443 7531
rect 23566 7528 23572 7540
rect 23431 7500 23572 7528
rect 23431 7497 23443 7500
rect 23385 7491 23443 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 25038 7488 25044 7540
rect 25096 7528 25102 7540
rect 26329 7531 26387 7537
rect 26329 7528 26341 7531
rect 25096 7500 26341 7528
rect 25096 7488 25102 7500
rect 26329 7497 26341 7500
rect 26375 7528 26387 7531
rect 26418 7528 26424 7540
rect 26375 7500 26424 7528
rect 26375 7497 26387 7500
rect 26329 7491 26387 7497
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 27157 7531 27215 7537
rect 27157 7497 27169 7531
rect 27203 7497 27215 7531
rect 27157 7491 27215 7497
rect 15841 7463 15899 7469
rect 15841 7429 15853 7463
rect 15887 7460 15899 7463
rect 16942 7460 16948 7472
rect 15887 7432 16948 7460
rect 15887 7429 15899 7432
rect 15841 7423 15899 7429
rect 16942 7420 16948 7432
rect 17000 7420 17006 7472
rect 17678 7420 17684 7472
rect 17736 7460 17742 7472
rect 17957 7463 18015 7469
rect 17957 7460 17969 7463
rect 17736 7432 17969 7460
rect 17736 7420 17742 7432
rect 17957 7429 17969 7432
rect 18003 7429 18015 7463
rect 17957 7423 18015 7429
rect 18173 7463 18231 7469
rect 18173 7429 18185 7463
rect 18219 7460 18231 7463
rect 18506 7460 18512 7472
rect 18219 7432 18512 7460
rect 18219 7429 18231 7432
rect 18173 7423 18231 7429
rect 18506 7420 18512 7432
rect 18564 7420 18570 7472
rect 20714 7460 20720 7472
rect 19996 7432 20720 7460
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 18966 7392 18972 7404
rect 16684 7364 18972 7392
rect 16684 7336 16712 7364
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19245 7395 19303 7401
rect 19245 7361 19257 7395
rect 19291 7361 19303 7395
rect 19426 7392 19432 7404
rect 19387 7364 19432 7392
rect 19245 7355 19303 7361
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 2774 7324 2780 7336
rect 2735 7296 2780 7324
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 16025 7327 16083 7333
rect 16025 7293 16037 7327
rect 16071 7293 16083 7327
rect 16666 7324 16672 7336
rect 16627 7296 16672 7324
rect 16025 7287 16083 7293
rect 16040 7256 16068 7287
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 16850 7256 16856 7268
rect 16040 7228 16856 7256
rect 16850 7216 16856 7228
rect 16908 7256 16914 7268
rect 16960 7256 16988 7287
rect 17034 7284 17040 7336
rect 17092 7324 17098 7336
rect 18506 7324 18512 7336
rect 17092 7296 18512 7324
rect 17092 7284 17098 7296
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 19260 7324 19288 7355
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 19518 7352 19524 7404
rect 19576 7392 19582 7404
rect 19996 7401 20024 7432
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 20898 7460 20904 7472
rect 20859 7432 20904 7460
rect 20898 7420 20904 7432
rect 20956 7420 20962 7472
rect 20993 7463 21051 7469
rect 20993 7429 21005 7463
rect 21039 7460 21051 7463
rect 21450 7460 21456 7472
rect 21039 7432 21456 7460
rect 21039 7429 21051 7432
rect 20993 7423 21051 7429
rect 21450 7420 21456 7432
rect 21508 7460 21514 7472
rect 22370 7460 22376 7472
rect 21508 7432 22376 7460
rect 21508 7420 21514 7432
rect 22370 7420 22376 7432
rect 22428 7420 22434 7472
rect 27172 7460 27200 7491
rect 27246 7488 27252 7540
rect 27304 7528 27310 7540
rect 28442 7528 28448 7540
rect 27304 7500 28448 7528
rect 27304 7488 27310 7500
rect 26344 7432 27200 7460
rect 26344 7404 26372 7432
rect 19981 7395 20039 7401
rect 19576 7364 19621 7392
rect 19576 7352 19582 7364
rect 19981 7361 19993 7395
rect 20027 7361 20039 7395
rect 20162 7392 20168 7404
rect 20123 7364 20168 7392
rect 19981 7355 20039 7361
rect 20162 7352 20168 7364
rect 20220 7352 20226 7404
rect 20806 7392 20812 7404
rect 20767 7364 20812 7392
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 21111 7395 21169 7401
rect 21111 7392 21123 7395
rect 21100 7361 21123 7392
rect 21157 7361 21169 7395
rect 22002 7392 22008 7404
rect 21963 7364 22008 7392
rect 21100 7355 21169 7361
rect 20346 7324 20352 7336
rect 19260 7296 20352 7324
rect 20346 7284 20352 7296
rect 20404 7284 20410 7336
rect 17678 7256 17684 7268
rect 16908 7228 17684 7256
rect 16908 7216 16914 7228
rect 17678 7216 17684 7228
rect 17736 7216 17742 7268
rect 18325 7259 18383 7265
rect 18325 7225 18337 7259
rect 18371 7256 18383 7259
rect 19334 7256 19340 7268
rect 18371 7228 19340 7256
rect 18371 7225 18383 7228
rect 18325 7219 18383 7225
rect 19334 7216 19340 7228
rect 19392 7216 19398 7268
rect 21100 7256 21128 7355
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7392 22891 7395
rect 23014 7392 23020 7404
rect 22879 7364 23020 7392
rect 22879 7361 22891 7364
rect 22833 7355 22891 7361
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 23198 7392 23204 7404
rect 23159 7364 23204 7392
rect 23198 7352 23204 7364
rect 23256 7352 23262 7404
rect 23290 7352 23296 7404
rect 23348 7392 23354 7404
rect 24029 7395 24087 7401
rect 24029 7392 24041 7395
rect 23348 7364 24041 7392
rect 23348 7352 23354 7364
rect 24029 7361 24041 7364
rect 24075 7361 24087 7395
rect 24029 7355 24087 7361
rect 24486 7352 24492 7404
rect 24544 7392 24550 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 24544 7364 24685 7392
rect 24544 7352 24550 7364
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 24949 7395 25007 7401
rect 24949 7392 24961 7395
rect 24912 7364 24961 7392
rect 24912 7352 24918 7364
rect 24949 7361 24961 7364
rect 24995 7361 25007 7395
rect 25130 7392 25136 7404
rect 25091 7364 25136 7392
rect 24949 7355 25007 7361
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 25774 7352 25780 7404
rect 25832 7392 25838 7404
rect 25961 7395 26019 7401
rect 25961 7392 25973 7395
rect 25832 7364 25973 7392
rect 25832 7352 25838 7364
rect 25961 7361 25973 7364
rect 26007 7361 26019 7395
rect 26142 7392 26148 7404
rect 26103 7364 26148 7392
rect 25961 7355 26019 7361
rect 26142 7352 26148 7364
rect 26200 7352 26206 7404
rect 26326 7352 26332 7404
rect 26384 7352 26390 7404
rect 27062 7352 27068 7404
rect 27120 7392 27126 7404
rect 27154 7395 27212 7401
rect 27154 7392 27166 7395
rect 27120 7364 27166 7392
rect 27120 7352 27126 7364
rect 27154 7361 27166 7364
rect 27200 7392 27212 7395
rect 27338 7392 27344 7404
rect 27200 7364 27344 7392
rect 27200 7361 27212 7364
rect 27154 7355 27212 7361
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 27448 7392 27476 7500
rect 28442 7488 28448 7500
rect 28500 7488 28506 7540
rect 27798 7420 27804 7472
rect 27856 7460 27862 7472
rect 28537 7463 28595 7469
rect 28537 7460 28549 7463
rect 27856 7432 28549 7460
rect 27856 7420 27862 7432
rect 28537 7429 28549 7432
rect 28583 7429 28595 7463
rect 28537 7423 28595 7429
rect 27617 7395 27675 7401
rect 27617 7392 27629 7395
rect 27448 7364 27629 7392
rect 27617 7361 27629 7364
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 29638 7352 29644 7404
rect 29696 7352 29702 7404
rect 35618 7392 35624 7404
rect 35579 7364 35624 7392
rect 35618 7352 35624 7364
rect 35676 7352 35682 7404
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21315 7296 21833 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21821 7293 21833 7296
rect 21867 7324 21879 7327
rect 22094 7324 22100 7336
rect 21867 7296 22100 7324
rect 21867 7293 21879 7296
rect 21821 7287 21879 7293
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 22738 7324 22744 7336
rect 22651 7296 22744 7324
rect 22738 7284 22744 7296
rect 22796 7324 22802 7336
rect 24118 7324 24124 7336
rect 22796 7296 24124 7324
rect 22796 7284 22802 7296
rect 24118 7284 24124 7296
rect 24176 7324 24182 7336
rect 27080 7324 27108 7352
rect 24176 7296 27108 7324
rect 24176 7284 24182 7296
rect 27430 7284 27436 7336
rect 27488 7324 27494 7336
rect 27525 7327 27583 7333
rect 27525 7324 27537 7327
rect 27488 7296 27537 7324
rect 27488 7284 27494 7296
rect 27525 7293 27537 7296
rect 27571 7293 27583 7327
rect 27525 7287 27583 7293
rect 27706 7284 27712 7336
rect 27764 7324 27770 7336
rect 28258 7324 28264 7336
rect 27764 7296 28264 7324
rect 27764 7284 27770 7296
rect 28258 7284 28264 7296
rect 28316 7284 28322 7336
rect 22922 7256 22928 7268
rect 21100 7228 22928 7256
rect 22922 7216 22928 7228
rect 22980 7216 22986 7268
rect 23842 7256 23848 7268
rect 23755 7228 23848 7256
rect 23842 7216 23848 7228
rect 23900 7256 23906 7268
rect 25314 7256 25320 7268
rect 23900 7228 25320 7256
rect 23900 7216 23906 7228
rect 25314 7216 25320 7228
rect 25372 7216 25378 7268
rect 15378 7188 15384 7200
rect 15339 7160 15384 7188
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 18141 7191 18199 7197
rect 18141 7157 18153 7191
rect 18187 7188 18199 7191
rect 18414 7188 18420 7200
rect 18187 7160 18420 7188
rect 18187 7157 18199 7160
rect 18141 7151 18199 7157
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 18506 7148 18512 7200
rect 18564 7188 18570 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18564 7160 19073 7188
rect 18564 7148 18570 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 20622 7188 20628 7200
rect 20583 7160 20628 7188
rect 19061 7151 19119 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 23198 7188 23204 7200
rect 23159 7160 23204 7188
rect 23198 7148 23204 7160
rect 23256 7148 23262 7200
rect 24762 7148 24768 7200
rect 24820 7197 24826 7200
rect 24820 7191 24869 7197
rect 24820 7157 24823 7191
rect 24857 7157 24869 7191
rect 24820 7151 24869 7157
rect 25041 7191 25099 7197
rect 25041 7157 25053 7191
rect 25087 7188 25099 7191
rect 26234 7188 26240 7200
rect 25087 7160 26240 7188
rect 25087 7157 25099 7160
rect 25041 7151 25099 7157
rect 24820 7148 24826 7151
rect 26234 7148 26240 7160
rect 26292 7148 26298 7200
rect 26970 7188 26976 7200
rect 26931 7160 26976 7188
rect 26970 7148 26976 7160
rect 27028 7148 27034 7200
rect 28994 7148 29000 7200
rect 29052 7188 29058 7200
rect 30009 7191 30067 7197
rect 30009 7188 30021 7191
rect 29052 7160 30021 7188
rect 29052 7148 29058 7160
rect 30009 7157 30021 7160
rect 30055 7157 30067 7191
rect 30009 7151 30067 7157
rect 36262 7148 36268 7200
rect 36320 7188 36326 7200
rect 37645 7191 37703 7197
rect 37645 7188 37657 7191
rect 36320 7160 37657 7188
rect 36320 7148 36326 7160
rect 37645 7157 37657 7160
rect 37691 7157 37703 7191
rect 37645 7151 37703 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2225 6987 2283 6993
rect 2225 6984 2237 6987
rect 2004 6956 2237 6984
rect 2004 6944 2010 6956
rect 2225 6953 2237 6956
rect 2271 6953 2283 6987
rect 2225 6947 2283 6953
rect 22465 6987 22523 6993
rect 22465 6953 22477 6987
rect 22511 6984 22523 6987
rect 22738 6984 22744 6996
rect 22511 6956 22744 6984
rect 22511 6953 22523 6956
rect 22465 6947 22523 6953
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 26786 6944 26792 6996
rect 26844 6984 26850 6996
rect 27890 6984 27896 6996
rect 26844 6956 27896 6984
rect 26844 6944 26850 6956
rect 27890 6944 27896 6956
rect 27948 6993 27954 6996
rect 27948 6987 27997 6993
rect 27948 6953 27951 6987
rect 27985 6953 27997 6987
rect 27948 6947 27997 6953
rect 27948 6944 27954 6947
rect 18601 6919 18659 6925
rect 18601 6885 18613 6919
rect 18647 6885 18659 6919
rect 18601 6879 18659 6885
rect 21913 6919 21971 6925
rect 21913 6885 21925 6919
rect 21959 6885 21971 6919
rect 21913 6879 21971 6885
rect 25332 6888 26924 6916
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6848 14611 6851
rect 15838 6848 15844 6860
rect 14599 6820 15844 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16666 6848 16672 6860
rect 16347 6820 16672 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 17034 6808 17040 6860
rect 17092 6848 17098 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 17092 6820 17141 6848
rect 17092 6808 17098 6820
rect 17129 6817 17141 6820
rect 17175 6848 17187 6851
rect 18230 6848 18236 6860
rect 17175 6820 18236 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 18616 6848 18644 6879
rect 20622 6848 20628 6860
rect 18616 6820 20628 6848
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 21266 6808 21272 6860
rect 21324 6848 21330 6860
rect 21928 6848 21956 6879
rect 21324 6820 21956 6848
rect 22281 6851 22339 6857
rect 21324 6808 21330 6820
rect 22281 6817 22293 6851
rect 22327 6848 22339 6851
rect 23198 6848 23204 6860
rect 22327 6820 23204 6848
rect 22327 6817 22339 6820
rect 22281 6811 22339 6817
rect 23198 6808 23204 6820
rect 23256 6848 23262 6860
rect 25332 6848 25360 6888
rect 25498 6848 25504 6860
rect 23256 6820 25360 6848
rect 25459 6820 25504 6848
rect 23256 6808 23262 6820
rect 25498 6808 25504 6820
rect 25556 6848 25562 6860
rect 26896 6848 26924 6888
rect 27709 6851 27767 6857
rect 27709 6848 27721 6851
rect 25556 6820 26832 6848
rect 26896 6820 27721 6848
rect 25556 6808 25562 6820
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6749 2375 6783
rect 2958 6780 2964 6792
rect 2919 6752 2964 6780
rect 2317 6743 2375 6749
rect 2332 6712 2360 6743
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 16942 6780 16948 6792
rect 16903 6752 16948 6780
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 18414 6780 18420 6792
rect 17267 6752 18420 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6749 19487 6783
rect 20898 6780 20904 6792
rect 20859 6752 20904 6780
rect 19429 6743 19487 6749
rect 5626 6712 5632 6724
rect 2332 6684 5632 6712
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 14826 6712 14832 6724
rect 14787 6684 14832 6712
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 15470 6672 15476 6724
rect 15528 6672 15534 6724
rect 19444 6712 19472 6743
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 21082 6780 21088 6792
rect 21043 6752 21088 6780
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6780 21419 6783
rect 21450 6780 21456 6792
rect 21407 6752 21456 6780
rect 21407 6749 21419 6752
rect 21361 6743 21419 6749
rect 21450 6740 21456 6752
rect 21508 6740 21514 6792
rect 22002 6740 22008 6792
rect 22060 6780 22066 6792
rect 22097 6783 22155 6789
rect 22097 6780 22109 6783
rect 22060 6752 22109 6780
rect 22060 6740 22066 6752
rect 22097 6749 22109 6752
rect 22143 6749 22155 6783
rect 22097 6743 22155 6749
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 22557 6783 22615 6789
rect 22557 6780 22569 6783
rect 22244 6752 22569 6780
rect 22244 6740 22250 6752
rect 22557 6749 22569 6752
rect 22603 6749 22615 6783
rect 22557 6743 22615 6749
rect 23017 6783 23075 6789
rect 23017 6749 23029 6783
rect 23063 6780 23075 6783
rect 23106 6780 23112 6792
rect 23063 6752 23112 6780
rect 23063 6749 23075 6752
rect 23017 6743 23075 6749
rect 23106 6740 23112 6752
rect 23164 6740 23170 6792
rect 23382 6780 23388 6792
rect 23295 6752 23388 6780
rect 23382 6740 23388 6752
rect 23440 6780 23446 6792
rect 24670 6780 24676 6792
rect 23440 6752 24676 6780
rect 23440 6740 23446 6752
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 25038 6740 25044 6792
rect 25096 6780 25102 6792
rect 25222 6780 25228 6792
rect 25096 6752 25228 6780
rect 25096 6740 25102 6752
rect 25222 6740 25228 6752
rect 25280 6780 25286 6792
rect 25409 6783 25467 6789
rect 25409 6780 25421 6783
rect 25280 6752 25421 6780
rect 25280 6740 25286 6752
rect 25409 6749 25421 6752
rect 25455 6780 25467 6783
rect 26145 6783 26203 6789
rect 26145 6780 26157 6783
rect 25455 6752 26157 6780
rect 25455 6749 25467 6752
rect 25409 6743 25467 6749
rect 26145 6749 26157 6752
rect 26191 6749 26203 6783
rect 26326 6780 26332 6792
rect 26287 6752 26332 6780
rect 26145 6743 26203 6749
rect 26326 6740 26332 6752
rect 26384 6740 26390 6792
rect 26804 6789 26832 6820
rect 27709 6817 27721 6820
rect 27755 6848 27767 6851
rect 28994 6848 29000 6860
rect 27755 6820 29000 6848
rect 27755 6817 27767 6820
rect 27709 6811 27767 6817
rect 28994 6808 29000 6820
rect 29052 6808 29058 6860
rect 29638 6848 29644 6860
rect 29599 6820 29644 6848
rect 29638 6808 29644 6820
rect 29696 6808 29702 6860
rect 36262 6848 36268 6860
rect 36223 6820 36268 6848
rect 36262 6808 36268 6820
rect 36320 6808 36326 6860
rect 37182 6848 37188 6860
rect 37143 6820 37188 6848
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6749 26847 6783
rect 26970 6780 26976 6792
rect 26931 6752 26976 6780
rect 26789 6743 26847 6749
rect 26970 6740 26976 6752
rect 27028 6740 27034 6792
rect 29733 6783 29791 6789
rect 29733 6749 29745 6783
rect 29779 6780 29791 6783
rect 30374 6780 30380 6792
rect 29779 6752 30380 6780
rect 29779 6749 29791 6752
rect 29733 6743 29791 6749
rect 30374 6740 30380 6752
rect 30432 6740 30438 6792
rect 19978 6712 19984 6724
rect 19444 6684 19984 6712
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 20990 6712 20996 6724
rect 20951 6684 20996 6712
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 21174 6672 21180 6724
rect 21232 6721 21238 6724
rect 21232 6715 21261 6721
rect 21249 6681 21261 6715
rect 23290 6712 23296 6724
rect 23251 6684 23296 6712
rect 21232 6675 21261 6681
rect 21232 6672 21238 6675
rect 23290 6672 23296 6684
rect 23348 6672 23354 6724
rect 25317 6715 25375 6721
rect 25317 6681 25329 6715
rect 25363 6712 25375 6715
rect 26237 6715 26295 6721
rect 26237 6712 26249 6715
rect 25363 6684 26249 6712
rect 25363 6681 25375 6684
rect 25317 6675 25375 6681
rect 26237 6681 26249 6684
rect 26283 6681 26295 6715
rect 36446 6712 36452 6724
rect 36407 6684 36452 6712
rect 26237 6675 26295 6681
rect 36446 6672 36452 6684
rect 36504 6672 36510 6724
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 1912 6616 2881 6644
rect 1912 6604 1918 6616
rect 2869 6613 2881 6616
rect 2915 6613 2927 6647
rect 16758 6644 16764 6656
rect 16719 6616 16764 6644
rect 2869 6607 2927 6613
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 18782 6604 18788 6656
rect 18840 6644 18846 6656
rect 19659 6647 19717 6653
rect 19659 6644 19671 6647
rect 18840 6616 19671 6644
rect 18840 6604 18846 6616
rect 19659 6613 19671 6616
rect 19705 6613 19717 6647
rect 19659 6607 19717 6613
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 20717 6647 20775 6653
rect 20717 6644 20729 6647
rect 20680 6616 20729 6644
rect 20680 6604 20686 6616
rect 20717 6613 20729 6616
rect 20763 6613 20775 6647
rect 20717 6607 20775 6613
rect 22462 6604 22468 6656
rect 22520 6644 22526 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22520 6616 23029 6644
rect 22520 6604 22526 6616
rect 23017 6613 23029 6616
rect 23063 6613 23075 6647
rect 23017 6607 23075 6613
rect 23106 6604 23112 6656
rect 23164 6644 23170 6656
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 23164 6616 23213 6644
rect 23164 6604 23170 6616
rect 23201 6613 23213 6616
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 24949 6647 25007 6653
rect 24949 6613 24961 6647
rect 24995 6644 25007 6647
rect 25222 6644 25228 6656
rect 24995 6616 25228 6644
rect 24995 6613 25007 6616
rect 24949 6607 25007 6613
rect 25222 6604 25228 6616
rect 25280 6604 25286 6656
rect 26881 6647 26939 6653
rect 26881 6613 26893 6647
rect 26927 6644 26939 6647
rect 28534 6644 28540 6656
rect 26927 6616 28540 6644
rect 26927 6613 26939 6616
rect 26881 6607 26939 6613
rect 28534 6604 28540 6616
rect 28592 6604 28598 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 14884 6412 15117 6440
rect 14884 6400 14890 6412
rect 15105 6409 15117 6412
rect 15151 6409 15163 6443
rect 15105 6403 15163 6409
rect 17034 6400 17040 6452
rect 17092 6449 17098 6452
rect 17092 6443 17111 6449
rect 17099 6409 17111 6443
rect 17092 6403 17111 6409
rect 17092 6400 17098 6403
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 20990 6440 20996 6452
rect 18012 6412 19012 6440
rect 20951 6412 20996 6440
rect 18012 6400 18018 6412
rect 1854 6372 1860 6384
rect 1815 6344 1860 6372
rect 1854 6332 1860 6344
rect 1912 6332 1918 6384
rect 16850 6372 16856 6384
rect 16811 6344 16856 6372
rect 16850 6332 16856 6344
rect 16908 6332 16914 6384
rect 18138 6372 18144 6384
rect 17972 6344 18144 6372
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15378 6304 15384 6316
rect 15335 6276 15384 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 17678 6304 17684 6316
rect 17236 6276 17684 6304
rect 2774 6236 2780 6248
rect 2735 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 17236 6177 17264 6276
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 17972 6313 18000 6344
rect 18138 6332 18144 6344
rect 18196 6372 18202 6384
rect 18782 6372 18788 6384
rect 18196 6344 18788 6372
rect 18196 6332 18202 6344
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 18984 6316 19012 6412
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 23566 6440 23572 6452
rect 22848 6412 23572 6440
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 20346 6372 20352 6384
rect 20036 6344 20352 6372
rect 20036 6332 20042 6344
rect 20346 6332 20352 6344
rect 20404 6372 20410 6384
rect 20441 6375 20499 6381
rect 20441 6372 20453 6375
rect 20404 6344 20453 6372
rect 20404 6332 20410 6344
rect 20441 6341 20453 6344
rect 20487 6341 20499 6375
rect 20441 6335 20499 6341
rect 20898 6332 20904 6384
rect 20956 6372 20962 6384
rect 22189 6375 22247 6381
rect 22189 6372 22201 6375
rect 20956 6344 22201 6372
rect 20956 6332 20962 6344
rect 22189 6341 22201 6344
rect 22235 6341 22247 6375
rect 22189 6335 22247 6341
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6273 17923 6307
rect 17865 6267 17923 6273
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 17880 6236 17908 6267
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18506 6304 18512 6316
rect 18104 6276 18512 6304
rect 18104 6264 18110 6276
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18966 6304 18972 6316
rect 18616 6276 18812 6304
rect 18879 6276 18972 6304
rect 18616 6236 18644 6276
rect 17880 6208 18644 6236
rect 18693 6239 18751 6245
rect 18693 6205 18705 6239
rect 18739 6205 18751 6239
rect 18784 6236 18812 6276
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 20993 6307 21051 6313
rect 20993 6273 21005 6307
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 18784 6208 19993 6236
rect 18693 6199 18751 6205
rect 19981 6205 19993 6208
rect 20027 6236 20039 6239
rect 20438 6236 20444 6248
rect 20027 6208 20444 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 17221 6171 17279 6177
rect 17221 6137 17233 6171
rect 17267 6137 17279 6171
rect 18414 6168 18420 6180
rect 17221 6131 17279 6137
rect 17512 6140 18420 6168
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 17037 6103 17095 6109
rect 17037 6100 17049 6103
rect 16724 6072 17049 6100
rect 16724 6060 16730 6072
rect 17037 6069 17049 6072
rect 17083 6100 17095 6103
rect 17512 6100 17540 6140
rect 18414 6128 18420 6140
rect 18472 6128 18478 6180
rect 18598 6128 18604 6180
rect 18656 6168 18662 6180
rect 18708 6168 18736 6199
rect 20438 6196 20444 6208
rect 20496 6196 20502 6248
rect 21008 6236 21036 6267
rect 21082 6264 21088 6316
rect 21140 6304 21146 6316
rect 22848 6313 22876 6412
rect 23566 6400 23572 6412
rect 23624 6440 23630 6452
rect 24026 6440 24032 6452
rect 23624 6412 24032 6440
rect 23624 6400 23630 6412
rect 24026 6400 24032 6412
rect 24084 6400 24090 6452
rect 25038 6440 25044 6452
rect 24999 6412 25044 6440
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 25130 6400 25136 6452
rect 25188 6440 25194 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 25188 6412 25513 6440
rect 25188 6400 25194 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 27062 6440 27068 6452
rect 27023 6412 27068 6440
rect 25501 6403 25559 6409
rect 27062 6400 27068 6412
rect 27120 6400 27126 6452
rect 23109 6375 23167 6381
rect 23109 6341 23121 6375
rect 23155 6372 23167 6375
rect 23934 6372 23940 6384
rect 23155 6344 23940 6372
rect 23155 6341 23167 6344
rect 23109 6335 23167 6341
rect 23934 6332 23940 6344
rect 23992 6372 23998 6384
rect 23992 6344 24164 6372
rect 23992 6332 23998 6344
rect 21177 6307 21235 6313
rect 21177 6304 21189 6307
rect 21140 6276 21189 6304
rect 21140 6264 21146 6276
rect 21177 6273 21189 6276
rect 21223 6304 21235 6307
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 21223 6276 21833 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 23017 6307 23075 6313
rect 23017 6273 23029 6307
rect 23063 6273 23075 6307
rect 23017 6267 23075 6273
rect 23201 6307 23259 6313
rect 23201 6273 23213 6307
rect 23247 6273 23259 6307
rect 23201 6267 23259 6273
rect 21450 6236 21456 6248
rect 21008 6208 21456 6236
rect 21450 6196 21456 6208
rect 21508 6236 21514 6248
rect 22020 6236 22048 6267
rect 21508 6208 22048 6236
rect 23032 6236 23060 6267
rect 23216 6236 23244 6267
rect 23750 6264 23756 6316
rect 23808 6304 23814 6316
rect 24136 6313 24164 6344
rect 27798 6332 27804 6384
rect 27856 6332 27862 6384
rect 28534 6372 28540 6384
rect 28495 6344 28540 6372
rect 28534 6332 28540 6344
rect 28592 6332 28598 6384
rect 37090 6332 37096 6384
rect 37148 6372 37154 6384
rect 37645 6375 37703 6381
rect 37645 6372 37657 6375
rect 37148 6344 37657 6372
rect 37148 6332 37154 6344
rect 37645 6341 37657 6344
rect 37691 6341 37703 6375
rect 37645 6335 37703 6341
rect 23845 6307 23903 6313
rect 23845 6304 23857 6307
rect 23808 6276 23857 6304
rect 23808 6264 23814 6276
rect 23845 6273 23857 6276
rect 23891 6273 23903 6307
rect 23845 6267 23903 6273
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6304 24179 6307
rect 24762 6304 24768 6316
rect 24167 6276 24768 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 24762 6264 24768 6276
rect 24820 6264 24826 6316
rect 24857 6307 24915 6313
rect 24857 6273 24869 6307
rect 24903 6273 24915 6307
rect 24857 6267 24915 6273
rect 23032 6208 23152 6236
rect 23216 6208 23888 6236
rect 21508 6196 21514 6208
rect 23124 6180 23152 6208
rect 19150 6168 19156 6180
rect 18656 6140 19156 6168
rect 18656 6128 18662 6140
rect 19150 6128 19156 6140
rect 19208 6168 19214 6180
rect 20073 6171 20131 6177
rect 20073 6168 20085 6171
rect 19208 6140 20085 6168
rect 19208 6128 19214 6140
rect 20073 6137 20085 6140
rect 20119 6137 20131 6171
rect 20073 6131 20131 6137
rect 23106 6128 23112 6180
rect 23164 6128 23170 6180
rect 23860 6112 23888 6208
rect 24670 6196 24676 6248
rect 24728 6236 24734 6248
rect 24872 6236 24900 6267
rect 25314 6264 25320 6316
rect 25372 6304 25378 6316
rect 25501 6307 25559 6313
rect 25501 6304 25513 6307
rect 25372 6276 25513 6304
rect 25372 6264 25378 6276
rect 25501 6273 25513 6276
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 25685 6307 25743 6313
rect 25685 6273 25697 6307
rect 25731 6304 25743 6307
rect 26510 6304 26516 6316
rect 25731 6276 26516 6304
rect 25731 6273 25743 6276
rect 25685 6267 25743 6273
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 28810 6264 28816 6316
rect 28868 6304 28874 6316
rect 38010 6304 38016 6316
rect 28868 6276 28913 6304
rect 37971 6276 38016 6304
rect 28868 6264 28874 6276
rect 38010 6264 38016 6276
rect 38068 6264 38074 6316
rect 24728 6208 24900 6236
rect 24728 6196 24734 6208
rect 17083 6072 17540 6100
rect 18233 6103 18291 6109
rect 17083 6069 17095 6072
rect 17037 6063 17095 6069
rect 18233 6069 18245 6103
rect 18279 6100 18291 6103
rect 19886 6100 19892 6112
rect 18279 6072 19892 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 19886 6060 19892 6072
rect 19944 6060 19950 6112
rect 23385 6103 23443 6109
rect 23385 6069 23397 6103
rect 23431 6100 23443 6103
rect 23474 6100 23480 6112
rect 23431 6072 23480 6100
rect 23431 6069 23443 6072
rect 23385 6063 23443 6069
rect 23474 6060 23480 6072
rect 23532 6060 23538 6112
rect 23842 6100 23848 6112
rect 23803 6072 23848 6100
rect 23842 6060 23848 6072
rect 23900 6060 23906 6112
rect 36722 6100 36728 6112
rect 36683 6072 36728 6100
rect 36722 6060 36728 6072
rect 36780 6060 36786 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 16666 5896 16672 5908
rect 16627 5868 16672 5896
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 17678 5896 17684 5908
rect 17639 5868 17684 5896
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 19426 5896 19432 5908
rect 19387 5868 19432 5896
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20312 5868 21680 5896
rect 20312 5856 20318 5868
rect 21652 5828 21680 5868
rect 22002 5856 22008 5908
rect 22060 5896 22066 5908
rect 22097 5899 22155 5905
rect 22097 5896 22109 5899
rect 22060 5868 22109 5896
rect 22060 5856 22066 5868
rect 22097 5865 22109 5868
rect 22143 5865 22155 5899
rect 22097 5859 22155 5865
rect 27709 5899 27767 5905
rect 27709 5865 27721 5899
rect 27755 5896 27767 5899
rect 27798 5896 27804 5908
rect 27755 5868 27804 5896
rect 27755 5865 27767 5868
rect 27709 5859 27767 5865
rect 27798 5856 27804 5868
rect 27856 5856 27862 5908
rect 21652 5800 24624 5828
rect 18046 5760 18052 5772
rect 17512 5732 18052 5760
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2038 5692 2044 5704
rect 1995 5664 2044 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2774 5692 2780 5704
rect 2639 5664 2780 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 3234 5692 3240 5704
rect 3195 5664 3240 5692
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 5040 5664 5089 5692
rect 5040 5652 5046 5664
rect 5077 5661 5089 5664
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 16022 5692 16028 5704
rect 15611 5664 16028 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16850 5692 16856 5704
rect 16811 5664 16856 5692
rect 16850 5652 16856 5664
rect 16908 5692 16914 5704
rect 17402 5692 17408 5704
rect 16908 5664 17408 5692
rect 16908 5652 16914 5664
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 17512 5701 17540 5732
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 18601 5763 18659 5769
rect 18601 5729 18613 5763
rect 18647 5760 18659 5763
rect 19334 5760 19340 5772
rect 18647 5732 19340 5760
rect 18647 5729 18659 5732
rect 18601 5723 18659 5729
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 20622 5760 20628 5772
rect 20583 5732 20628 5760
rect 20622 5720 20628 5732
rect 20680 5720 20686 5772
rect 23293 5763 23351 5769
rect 23293 5729 23305 5763
rect 23339 5760 23351 5763
rect 23566 5760 23572 5772
rect 23339 5732 23572 5760
rect 23339 5729 23351 5732
rect 23293 5723 23351 5729
rect 23566 5720 23572 5732
rect 23624 5720 23630 5772
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5692 17831 5695
rect 17954 5692 17960 5704
rect 17819 5664 17960 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 17954 5652 17960 5664
rect 18012 5652 18018 5704
rect 18506 5692 18512 5704
rect 18467 5664 18512 5692
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 18966 5652 18972 5704
rect 19024 5692 19030 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 19024 5664 19257 5692
rect 19024 5652 19030 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 19484 5664 20361 5692
rect 19484 5652 19490 5664
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 23014 5692 23020 5704
rect 22975 5664 23020 5692
rect 20349 5655 20407 5661
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 23842 5652 23848 5704
rect 23900 5692 23906 5704
rect 24596 5701 24624 5800
rect 37090 5760 37096 5772
rect 37051 5732 37096 5760
rect 37090 5720 37096 5732
rect 37148 5720 37154 5772
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 23900 5664 24409 5692
rect 23900 5652 23906 5664
rect 24397 5661 24409 5664
rect 24443 5661 24455 5695
rect 24397 5655 24455 5661
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 25222 5692 25228 5704
rect 25183 5664 25228 5692
rect 24581 5655 24639 5661
rect 25222 5652 25228 5664
rect 25280 5652 25286 5704
rect 25774 5652 25780 5704
rect 25832 5692 25838 5704
rect 25869 5695 25927 5701
rect 25869 5692 25881 5695
rect 25832 5664 25881 5692
rect 25832 5652 25838 5664
rect 25869 5661 25881 5664
rect 25915 5661 25927 5695
rect 25869 5655 25927 5661
rect 27801 5695 27859 5701
rect 27801 5661 27813 5695
rect 27847 5692 27859 5695
rect 30374 5692 30380 5704
rect 27847 5664 30380 5692
rect 27847 5661 27859 5664
rect 27801 5655 27859 5661
rect 30374 5652 30380 5664
rect 30432 5652 30438 5704
rect 34514 5652 34520 5704
rect 34572 5692 34578 5704
rect 35621 5695 35679 5701
rect 35621 5692 35633 5695
rect 34572 5664 35633 5692
rect 34572 5652 34578 5664
rect 35621 5661 35633 5664
rect 35667 5661 35679 5695
rect 35621 5655 35679 5661
rect 38102 5652 38108 5704
rect 38160 5692 38166 5704
rect 38160 5664 38205 5692
rect 38160 5652 38166 5664
rect 1857 5627 1915 5633
rect 1857 5593 1869 5627
rect 1903 5624 1915 5627
rect 3418 5624 3424 5636
rect 1903 5596 3424 5624
rect 1903 5593 1915 5596
rect 1857 5587 1915 5593
rect 3418 5584 3424 5596
rect 3476 5584 3482 5636
rect 19337 5627 19395 5633
rect 19337 5593 19349 5627
rect 19383 5593 19395 5627
rect 19337 5587 19395 5593
rect 19521 5627 19579 5633
rect 19521 5593 19533 5627
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 3050 5556 3056 5568
rect 2547 5528 3056 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 16117 5559 16175 5565
rect 16117 5525 16129 5559
rect 16163 5556 16175 5559
rect 16574 5556 16580 5568
rect 16163 5528 16580 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 17126 5516 17132 5568
rect 17184 5556 17190 5568
rect 17313 5559 17371 5565
rect 17313 5556 17325 5559
rect 17184 5528 17325 5556
rect 17184 5516 17190 5528
rect 17313 5525 17325 5528
rect 17359 5525 17371 5559
rect 17313 5519 17371 5525
rect 19242 5516 19248 5568
rect 19300 5556 19306 5568
rect 19352 5556 19380 5587
rect 19300 5528 19380 5556
rect 19536 5556 19564 5587
rect 20070 5584 20076 5636
rect 20128 5624 20134 5636
rect 37918 5624 37924 5636
rect 20128 5596 21114 5624
rect 37879 5596 37924 5624
rect 20128 5584 20134 5596
rect 37918 5584 37924 5596
rect 37976 5584 37982 5636
rect 20806 5556 20812 5568
rect 19536 5528 20812 5556
rect 19300 5516 19306 5528
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 23106 5516 23112 5568
rect 23164 5556 23170 5568
rect 24765 5559 24823 5565
rect 24765 5556 24777 5559
rect 23164 5528 24777 5556
rect 23164 5516 23170 5528
rect 24765 5525 24777 5528
rect 24811 5525 24823 5559
rect 24765 5519 24823 5525
rect 25317 5559 25375 5565
rect 25317 5525 25329 5559
rect 25363 5556 25375 5559
rect 25866 5556 25872 5568
rect 25363 5528 25872 5556
rect 25363 5525 25375 5528
rect 25317 5519 25375 5525
rect 25866 5516 25872 5528
rect 25924 5516 25930 5568
rect 25958 5516 25964 5568
rect 26016 5556 26022 5568
rect 26016 5528 26061 5556
rect 26016 5516 26022 5528
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 15933 5355 15991 5361
rect 15933 5321 15945 5355
rect 15979 5352 15991 5355
rect 16022 5352 16028 5364
rect 15979 5324 16028 5352
rect 15979 5321 15991 5324
rect 15933 5315 15991 5321
rect 16022 5312 16028 5324
rect 16080 5352 16086 5364
rect 18506 5352 18512 5364
rect 16080 5324 18512 5352
rect 16080 5312 16086 5324
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 18598 5312 18604 5364
rect 18656 5352 18662 5364
rect 18656 5324 18701 5352
rect 18656 5312 18662 5324
rect 20346 5312 20352 5364
rect 20404 5352 20410 5364
rect 23934 5361 23940 5364
rect 20809 5355 20867 5361
rect 20809 5352 20821 5355
rect 20404 5324 20821 5352
rect 20404 5312 20410 5324
rect 20809 5321 20821 5324
rect 20855 5321 20867 5355
rect 20809 5315 20867 5321
rect 22925 5355 22983 5361
rect 22925 5321 22937 5355
rect 22971 5352 22983 5355
rect 23753 5355 23811 5361
rect 23753 5352 23765 5355
rect 22971 5324 23765 5352
rect 22971 5321 22983 5324
rect 22925 5315 22983 5321
rect 23753 5321 23765 5324
rect 23799 5321 23811 5355
rect 23753 5315 23811 5321
rect 23921 5355 23940 5361
rect 23921 5321 23933 5355
rect 23921 5315 23940 5321
rect 23934 5312 23940 5315
rect 23992 5312 23998 5364
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 36446 5312 36452 5364
rect 36504 5352 36510 5364
rect 36633 5355 36691 5361
rect 36633 5352 36645 5355
rect 36504 5324 36645 5352
rect 36504 5312 36510 5324
rect 36633 5321 36645 5324
rect 36679 5321 36691 5355
rect 36633 5315 36691 5321
rect 37553 5355 37611 5361
rect 37553 5321 37565 5355
rect 37599 5352 37611 5355
rect 37918 5352 37924 5364
rect 37599 5324 37924 5352
rect 37599 5321 37611 5324
rect 37553 5315 37611 5321
rect 37918 5312 37924 5324
rect 37976 5312 37982 5364
rect 3418 5284 3424 5296
rect 3379 5256 3424 5284
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 17126 5284 17132 5296
rect 17087 5256 17132 5284
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 17862 5244 17868 5296
rect 17920 5244 17926 5296
rect 19334 5244 19340 5296
rect 19392 5284 19398 5296
rect 23017 5287 23075 5293
rect 19392 5256 19826 5284
rect 19392 5244 19398 5256
rect 23017 5253 23029 5287
rect 23063 5284 23075 5287
rect 23106 5284 23112 5296
rect 23063 5256 23112 5284
rect 23063 5253 23075 5256
rect 23017 5247 23075 5253
rect 23106 5244 23112 5256
rect 23164 5244 23170 5296
rect 23566 5244 23572 5296
rect 23624 5284 23630 5296
rect 24121 5287 24179 5293
rect 24121 5284 24133 5287
rect 23624 5256 24133 5284
rect 23624 5244 23630 5256
rect 24121 5253 24133 5256
rect 24167 5253 24179 5287
rect 24121 5247 24179 5253
rect 25682 5244 25688 5296
rect 25740 5244 25746 5296
rect 25866 5244 25872 5296
rect 25924 5284 25930 5296
rect 26145 5287 26203 5293
rect 26145 5284 26157 5287
rect 25924 5256 26157 5284
rect 25924 5244 25930 5256
rect 26145 5253 26157 5256
rect 26191 5253 26203 5287
rect 26145 5247 26203 5253
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3786 5216 3792 5228
rect 3651 5188 3792 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 5350 5216 5356 5228
rect 5311 5188 5356 5216
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 16114 5216 16120 5228
rect 16075 5188 16120 5216
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5185 22155 5219
rect 22097 5179 22155 5185
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 15930 5108 15936 5160
rect 15988 5148 15994 5160
rect 16853 5151 16911 5157
rect 16853 5148 16865 5151
rect 15988 5120 16865 5148
rect 15988 5108 15994 5120
rect 16853 5117 16865 5120
rect 16899 5117 16911 5151
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 16853 5111 16911 5117
rect 18156 5120 19073 5148
rect 4062 5012 4068 5024
rect 4023 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 5224 4984 5273 5012
rect 5224 4972 5230 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 5261 4975 5319 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 16868 5012 16896 5111
rect 18156 5012 18184 5120
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 19337 5151 19395 5157
rect 19337 5117 19349 5151
rect 19383 5148 19395 5151
rect 19978 5148 19984 5160
rect 19383 5120 19984 5148
rect 19383 5117 19395 5120
rect 19337 5111 19395 5117
rect 16868 4984 18184 5012
rect 19076 5012 19104 5111
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 20346 5040 20352 5092
rect 20404 5080 20410 5092
rect 22112 5080 22140 5179
rect 36630 5176 36636 5228
rect 36688 5216 36694 5228
rect 36725 5219 36783 5225
rect 36725 5216 36737 5219
rect 36688 5188 36737 5216
rect 36688 5176 36694 5188
rect 36725 5185 36737 5188
rect 36771 5216 36783 5219
rect 37461 5219 37519 5225
rect 37461 5216 37473 5219
rect 36771 5188 37473 5216
rect 36771 5185 36783 5188
rect 36725 5179 36783 5185
rect 37461 5185 37473 5188
rect 37507 5185 37519 5219
rect 37461 5179 37519 5185
rect 23198 5148 23204 5160
rect 23159 5120 23204 5148
rect 23198 5108 23204 5120
rect 23256 5108 23262 5160
rect 26418 5148 26424 5160
rect 26379 5120 26424 5148
rect 26418 5108 26424 5120
rect 26476 5148 26482 5160
rect 28258 5148 28264 5160
rect 26476 5120 28264 5148
rect 26476 5108 26482 5120
rect 28258 5108 28264 5120
rect 28316 5108 28322 5160
rect 20404 5052 22140 5080
rect 20404 5040 20410 5052
rect 19426 5012 19432 5024
rect 19076 4984 19432 5012
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 21913 5015 21971 5021
rect 21913 4981 21925 5015
rect 21959 5012 21971 5015
rect 22186 5012 22192 5024
rect 21959 4984 22192 5012
rect 21959 4981 21971 4984
rect 21913 4975 21971 4981
rect 22186 4972 22192 4984
rect 22244 4972 22250 5024
rect 22370 4972 22376 5024
rect 22428 5012 22434 5024
rect 22557 5015 22615 5021
rect 22557 5012 22569 5015
rect 22428 4984 22569 5012
rect 22428 4972 22434 4984
rect 22557 4981 22569 4984
rect 22603 4981 22615 5015
rect 22557 4975 22615 4981
rect 23658 4972 23664 5024
rect 23716 5012 23722 5024
rect 23937 5015 23995 5021
rect 23937 5012 23949 5015
rect 23716 4984 23949 5012
rect 23716 4972 23722 4984
rect 23937 4981 23949 4984
rect 23983 4981 23995 5015
rect 23937 4975 23995 4981
rect 32582 4972 32588 5024
rect 32640 5012 32646 5024
rect 32953 5015 33011 5021
rect 32953 5012 32965 5015
rect 32640 4984 32965 5012
rect 32640 4972 32646 4984
rect 32953 4981 32965 4984
rect 32999 4981 33011 5015
rect 32953 4975 33011 4981
rect 34790 4972 34796 5024
rect 34848 5012 34854 5024
rect 34977 5015 35035 5021
rect 34977 5012 34989 5015
rect 34848 4984 34989 5012
rect 34848 4972 34854 4984
rect 34977 4981 34989 4984
rect 35023 4981 35035 5015
rect 34977 4975 35035 4981
rect 36081 5015 36139 5021
rect 36081 4981 36093 5015
rect 36127 5012 36139 5015
rect 36630 5012 36636 5024
rect 36127 4984 36636 5012
rect 36127 4981 36139 4984
rect 36081 4975 36139 4981
rect 36630 4972 36636 4984
rect 36688 4972 36694 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 15552 4811 15610 4817
rect 15552 4777 15564 4811
rect 15598 4808 15610 4811
rect 16758 4808 16764 4820
rect 15598 4780 16764 4808
rect 15598 4777 15610 4780
rect 15552 4771 15610 4777
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 16850 4768 16856 4820
rect 16908 4808 16914 4820
rect 17037 4811 17095 4817
rect 17037 4808 17049 4811
rect 16908 4780 17049 4808
rect 16908 4768 16914 4780
rect 17037 4777 17049 4780
rect 17083 4777 17095 4811
rect 17862 4808 17868 4820
rect 17823 4780 17868 4808
rect 17037 4771 17095 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 20346 4808 20352 4820
rect 17972 4780 20352 4808
rect 6886 4712 12434 4740
rect 3050 4672 3056 4684
rect 3011 4644 3056 4672
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3234 4672 3240 4684
rect 3195 4644 3240 4672
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 4982 4672 4988 4684
rect 4943 4644 4988 4672
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5810 4672 5816 4684
rect 5771 4644 5816 4672
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 658 4496 664 4548
rect 716 4536 722 4548
rect 1397 4539 1455 4545
rect 1397 4536 1409 4539
rect 716 4508 1409 4536
rect 716 4496 722 4508
rect 1397 4505 1409 4508
rect 1443 4505 1455 4539
rect 1397 4499 1455 4505
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 3988 4536 4016 4567
rect 6886 4536 6914 4712
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10778 4672 10784 4684
rect 9999 4644 10784 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 7466 4604 7472 4616
rect 7427 4576 7472 4604
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 8938 4604 8944 4616
rect 8343 4576 8944 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 9088 4576 9137 4604
rect 9088 4564 9094 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 9125 4567 9183 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 2832 4508 6914 4536
rect 2832 4496 2838 4508
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4154 4468 4160 4480
rect 3927 4440 4160 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 10597 4471 10655 4477
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 11422 4468 11428 4480
rect 10643 4440 11428 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 12406 4468 12434 4712
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15930 4672 15936 4684
rect 15335 4644 15936 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 17972 4672 18000 4780
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 21177 4811 21235 4817
rect 21177 4777 21189 4811
rect 21223 4808 21235 4811
rect 22094 4808 22100 4820
rect 21223 4780 22100 4808
rect 21223 4777 21235 4780
rect 21177 4771 21235 4777
rect 22094 4768 22100 4780
rect 22152 4768 22158 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 23569 4811 23627 4817
rect 23569 4808 23581 4811
rect 23256 4780 23581 4808
rect 23256 4768 23262 4780
rect 23569 4777 23581 4780
rect 23615 4777 23627 4811
rect 23569 4771 23627 4777
rect 16172 4644 18000 4672
rect 18616 4712 19564 4740
rect 16172 4632 16178 4644
rect 17773 4607 17831 4613
rect 17773 4573 17785 4607
rect 17819 4604 17831 4607
rect 18506 4604 18512 4616
rect 17819 4576 18512 4604
rect 17819 4573 17831 4576
rect 17773 4567 17831 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 16574 4496 16580 4548
rect 16632 4496 16638 4548
rect 18616 4536 18644 4712
rect 19426 4672 19432 4684
rect 19387 4644 19432 4672
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 19536 4672 19564 4712
rect 23290 4700 23296 4752
rect 23348 4740 23354 4752
rect 25041 4743 25099 4749
rect 25041 4740 25053 4743
rect 23348 4712 25053 4740
rect 23348 4700 23354 4712
rect 25041 4709 25053 4712
rect 25087 4709 25099 4743
rect 25041 4703 25099 4709
rect 21726 4672 21732 4684
rect 19536 4644 21732 4672
rect 21726 4632 21732 4644
rect 21784 4632 21790 4684
rect 21821 4675 21879 4681
rect 21821 4641 21833 4675
rect 21867 4672 21879 4675
rect 24762 4672 24768 4684
rect 21867 4644 24768 4672
rect 21867 4641 21879 4644
rect 21821 4635 21879 4641
rect 24762 4632 24768 4644
rect 24820 4672 24826 4684
rect 26418 4672 26424 4684
rect 24820 4644 26424 4672
rect 24820 4632 24826 4644
rect 26418 4632 26424 4644
rect 26476 4672 26482 4684
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 26476 4644 26801 4672
rect 26476 4632 26482 4644
rect 26789 4641 26801 4644
rect 26835 4641 26847 4675
rect 33134 4672 33140 4684
rect 33095 4644 33140 4672
rect 26789 4635 26847 4641
rect 33134 4632 33140 4644
rect 33192 4632 33198 4684
rect 35713 4675 35771 4681
rect 35713 4641 35725 4675
rect 35759 4672 35771 4675
rect 37274 4672 37280 4684
rect 35759 4644 37280 4672
rect 35759 4641 35771 4644
rect 35713 4635 35771 4641
rect 37274 4632 37280 4644
rect 37332 4632 37338 4684
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 23440 4576 24593 4604
rect 23440 4564 23446 4576
rect 24581 4573 24593 4576
rect 24627 4604 24639 4607
rect 24627 4576 25176 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 16868 4508 18644 4536
rect 19705 4539 19763 4545
rect 16868 4468 16896 4508
rect 19705 4505 19717 4539
rect 19751 4536 19763 4539
rect 19978 4536 19984 4548
rect 19751 4508 19984 4536
rect 19751 4505 19763 4508
rect 19705 4499 19763 4505
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 20088 4508 20194 4536
rect 12406 4440 16896 4468
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 20088 4468 20116 4508
rect 22094 4496 22100 4548
rect 22152 4536 22158 4548
rect 22152 4508 22197 4536
rect 22152 4496 22158 4508
rect 23106 4496 23112 4548
rect 23164 4496 23170 4548
rect 24486 4468 24492 4480
rect 18647 4440 20116 4468
rect 24447 4440 24492 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 24486 4428 24492 4440
rect 24544 4428 24550 4480
rect 25148 4468 25176 4576
rect 31754 4564 31760 4616
rect 31812 4604 31818 4616
rect 32217 4607 32275 4613
rect 32217 4604 32229 4607
rect 31812 4576 32229 4604
rect 31812 4564 31818 4576
rect 32217 4573 32229 4576
rect 32263 4573 32275 4607
rect 32217 4567 32275 4573
rect 34698 4564 34704 4616
rect 34756 4604 34762 4616
rect 35069 4607 35127 4613
rect 35069 4604 35081 4607
rect 34756 4576 35081 4604
rect 34756 4564 34762 4576
rect 35069 4573 35081 4576
rect 35115 4573 35127 4607
rect 35069 4567 35127 4573
rect 25958 4496 25964 4548
rect 26016 4496 26022 4548
rect 26234 4496 26240 4548
rect 26292 4536 26298 4548
rect 26513 4539 26571 4545
rect 26513 4536 26525 4539
rect 26292 4508 26525 4536
rect 26292 4496 26298 4508
rect 26513 4505 26525 4508
rect 26559 4505 26571 4539
rect 32398 4536 32404 4548
rect 32359 4508 32404 4536
rect 26513 4499 26571 4505
rect 32398 4496 32404 4508
rect 32456 4496 32462 4548
rect 35161 4539 35219 4545
rect 35161 4505 35173 4539
rect 35207 4536 35219 4539
rect 35897 4539 35955 4545
rect 35897 4536 35909 4539
rect 35207 4508 35909 4536
rect 35207 4505 35219 4508
rect 35161 4499 35219 4505
rect 35897 4505 35909 4508
rect 35943 4505 35955 4539
rect 37550 4536 37556 4548
rect 37511 4508 37556 4536
rect 35897 4499 35955 4505
rect 37550 4496 37556 4508
rect 37608 4496 37614 4548
rect 25774 4468 25780 4480
rect 25148 4440 25780 4468
rect 25774 4428 25780 4440
rect 25832 4428 25838 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 19889 4267 19947 4273
rect 19889 4233 19901 4267
rect 19935 4264 19947 4267
rect 19978 4264 19984 4276
rect 19935 4236 19984 4264
rect 19935 4233 19947 4236
rect 19889 4227 19947 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 22189 4267 22247 4273
rect 22189 4264 22201 4267
rect 22152 4236 22201 4264
rect 22152 4224 22158 4236
rect 22189 4233 22201 4236
rect 22235 4233 22247 4267
rect 22189 4227 22247 4233
rect 3418 4156 3424 4208
rect 3476 4196 3482 4208
rect 24486 4196 24492 4208
rect 3476 4168 8892 4196
rect 3476 4156 3482 4168
rect 5166 4128 5172 4140
rect 5127 4100 5172 4128
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 4154 4060 4160 4072
rect 4115 4032 4160 4060
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8294 4060 8300 4072
rect 7699 4032 8300 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 4356 3992 4384 4023
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8864 4069 8892 4168
rect 19352 4168 19564 4196
rect 24058 4168 24492 4196
rect 9950 4128 9956 4140
rect 9911 4100 9956 4128
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10870 4128 10876 4140
rect 10643 4100 10876 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 19352 4128 19380 4168
rect 18748 4100 19380 4128
rect 19429 4131 19487 4137
rect 18748 4088 18754 4100
rect 19429 4097 19441 4131
rect 19475 4097 19487 4131
rect 19536 4128 19564 4168
rect 24486 4156 24492 4168
rect 24544 4156 24550 4208
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19536 4100 20085 4128
rect 19429 4091 19487 4097
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20714 4128 20720 4140
rect 20675 4100 20720 4128
rect 20073 4091 20131 4097
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4029 8907 4063
rect 19444 4060 19472 4091
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 22370 4128 22376 4140
rect 22331 4100 22376 4128
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 23198 4128 23204 4140
rect 22848 4100 23204 4128
rect 22186 4060 22192 4072
rect 19444 4032 22192 4060
rect 8849 4023 8907 4029
rect 22186 4020 22192 4032
rect 22244 4060 22250 4072
rect 22848 4060 22876 4100
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 24762 4088 24768 4140
rect 24820 4128 24826 4140
rect 25682 4128 25688 4140
rect 24820 4100 24865 4128
rect 25643 4100 25688 4128
rect 24820 4088 24826 4100
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 25774 4088 25780 4140
rect 25832 4128 25838 4140
rect 31021 4131 31079 4137
rect 25832 4100 25877 4128
rect 25832 4088 25838 4100
rect 31021 4097 31033 4131
rect 31067 4097 31079 4131
rect 32582 4128 32588 4140
rect 32543 4100 32588 4128
rect 31021 4091 31079 4097
rect 23014 4060 23020 4072
rect 22244 4032 22876 4060
rect 22975 4032 23020 4060
rect 22244 4020 22250 4032
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 23474 4020 23480 4072
rect 23532 4060 23538 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 23532 4032 24501 4060
rect 23532 4020 23538 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 2087 3964 4384 3992
rect 5077 3995 5135 4001
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 5077 3961 5089 3995
rect 5123 3992 5135 3995
rect 6546 3992 6552 4004
rect 5123 3964 6552 3992
rect 5123 3961 5135 3964
rect 5077 3955 5135 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 19337 3995 19395 4001
rect 19337 3961 19349 3995
rect 19383 3992 19395 3995
rect 20070 3992 20076 4004
rect 19383 3964 20076 3992
rect 19383 3961 19395 3964
rect 19337 3955 19395 3961
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 21634 3952 21640 4004
rect 21692 3992 21698 4004
rect 21692 3964 23520 3992
rect 21692 3952 21698 3964
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 5902 3924 5908 3936
rect 5859 3896 5908 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6328 3896 6377 3924
rect 6328 3884 6334 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9272 3896 9873 3924
rect 9272 3884 9278 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10594 3924 10600 3936
rect 10551 3896 10600 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11296 3896 11529 3924
rect 11296 3884 11302 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 13265 3927 13323 3933
rect 13265 3893 13277 3927
rect 13311 3924 13323 3927
rect 13814 3924 13820 3936
rect 13311 3896 13820 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 20809 3927 20867 3933
rect 20809 3893 20821 3927
rect 20855 3924 20867 3927
rect 22370 3924 22376 3936
rect 20855 3896 22376 3924
rect 20855 3893 20867 3896
rect 20809 3887 20867 3893
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 23492 3924 23520 3964
rect 31036 3924 31064 4091
rect 32582 4088 32588 4100
rect 32640 4088 32646 4140
rect 36722 4088 36728 4140
rect 36780 4128 36786 4140
rect 37274 4128 37280 4140
rect 36780 4100 36825 4128
rect 37235 4100 37280 4128
rect 36780 4088 36786 4100
rect 37274 4088 37280 4100
rect 37332 4088 37338 4140
rect 38102 4128 38108 4140
rect 38063 4100 38108 4128
rect 38102 4088 38108 4100
rect 38160 4088 38166 4140
rect 32769 4063 32827 4069
rect 32769 4029 32781 4063
rect 32815 4060 32827 4063
rect 33410 4060 33416 4072
rect 32815 4032 33416 4060
rect 32815 4029 32827 4032
rect 32769 4023 32827 4029
rect 33410 4020 33416 4032
rect 33468 4020 33474 4072
rect 33502 4020 33508 4072
rect 33560 4060 33566 4072
rect 35802 4060 35808 4072
rect 33560 4032 33605 4060
rect 35763 4032 35808 4060
rect 33560 4020 33566 4032
rect 35802 4020 35808 4032
rect 35860 4020 35866 4072
rect 36541 4063 36599 4069
rect 36541 4029 36553 4063
rect 36587 4060 36599 4063
rect 37826 4060 37832 4072
rect 36587 4032 37832 4060
rect 36587 4029 36599 4032
rect 36541 4023 36599 4029
rect 37826 4020 37832 4032
rect 37884 4020 37890 4072
rect 23492 3896 31064 3924
rect 31113 3927 31171 3933
rect 31113 3893 31125 3927
rect 31159 3924 31171 3927
rect 31202 3924 31208 3936
rect 31159 3896 31208 3924
rect 31159 3893 31171 3896
rect 31113 3887 31171 3893
rect 31202 3884 31208 3896
rect 31260 3884 31266 3936
rect 33594 3884 33600 3936
rect 33652 3924 33658 3936
rect 37918 3924 37924 3936
rect 33652 3896 37924 3924
rect 33652 3884 33658 3896
rect 37918 3884 37924 3896
rect 37976 3884 37982 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 8294 3720 8300 3732
rect 8255 3692 8300 3720
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 13354 3720 13360 3732
rect 8444 3692 13360 3720
rect 8444 3680 8450 3692
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 23106 3720 23112 3732
rect 23067 3692 23112 3720
rect 23106 3680 23112 3692
rect 23164 3680 23170 3732
rect 33410 3720 33416 3732
rect 33371 3692 33416 3720
rect 33410 3680 33416 3692
rect 33468 3680 33474 3732
rect 37826 3720 37832 3732
rect 37787 3692 37832 3720
rect 37826 3680 37832 3692
rect 37884 3680 37890 3732
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 3476 3624 8984 3652
rect 3476 3612 3482 3624
rect 4706 3584 4712 3596
rect 4667 3556 4712 3584
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 8956 3593 8984 3624
rect 10962 3612 10968 3664
rect 11020 3652 11026 3664
rect 32490 3652 32496 3664
rect 11020 3624 11744 3652
rect 11020 3612 11026 3624
rect 8941 3587 8999 3593
rect 6144 3556 8892 3584
rect 6144 3544 6150 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1762 3516 1768 3528
rect 1719 3488 1768 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 2958 3516 2964 3528
rect 2823 3488 2964 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 2332 3448 2360 3479
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 6052 3488 6377 3516
rect 6052 3476 6058 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 6365 3479 6423 3485
rect 6886 3488 7573 3516
rect 4154 3448 4160 3460
rect 2332 3420 4160 3448
rect 4154 3408 4160 3420
rect 4212 3408 4218 3460
rect 4338 3408 4344 3460
rect 4396 3448 4402 3460
rect 5721 3451 5779 3457
rect 5721 3448 5733 3451
rect 4396 3420 5733 3448
rect 4396 3408 4402 3420
rect 5721 3417 5733 3420
rect 5767 3417 5779 3451
rect 5721 3411 5779 3417
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2004 3352 2237 3380
rect 2004 3340 2010 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3380 2927 3383
rect 3050 3380 3056 3392
rect 2915 3352 3056 3380
rect 2915 3349 2927 3352
rect 2869 3343 2927 3349
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 6886 3380 6914 3488
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 8386 3516 8392 3528
rect 8347 3488 8392 3516
rect 7561 3479 7619 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 8864 3448 8892 3556
rect 8941 3553 8953 3587
rect 8987 3553 8999 3587
rect 10594 3584 10600 3596
rect 10555 3556 10600 3584
rect 8941 3547 8999 3553
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 10778 3584 10784 3596
rect 10739 3556 10784 3584
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11422 3584 11428 3596
rect 11383 3556 11428 3584
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 11716 3593 11744 3624
rect 19720 3624 32496 3652
rect 11701 3587 11759 3593
rect 11701 3553 11713 3587
rect 11747 3553 11759 3587
rect 11701 3547 11759 3553
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 15105 3587 15163 3593
rect 15105 3584 15117 3587
rect 14332 3556 15117 3584
rect 14332 3544 14338 3556
rect 15105 3553 15117 3556
rect 15151 3553 15163 3587
rect 15105 3547 15163 3553
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14608 3488 14657 3516
rect 14608 3476 14614 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 16298 3516 16304 3528
rect 16259 3488 16304 3516
rect 14645 3479 14703 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18966 3516 18972 3528
rect 18463 3488 18972 3516
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 17604 3448 17632 3479
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 19720 3525 19748 3624
rect 32490 3612 32496 3624
rect 32548 3612 32554 3664
rect 37918 3652 37924 3664
rect 35866 3624 37924 3652
rect 21174 3584 21180 3596
rect 21135 3556 21180 3584
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 22370 3584 22376 3596
rect 22331 3556 22376 3584
rect 22370 3544 22376 3556
rect 22428 3544 22434 3596
rect 31202 3584 31208 3596
rect 31163 3556 31208 3584
rect 31202 3544 31208 3556
rect 31260 3544 31266 3596
rect 31570 3584 31576 3596
rect 31531 3556 31576 3584
rect 31570 3544 31576 3556
rect 31628 3544 31634 3596
rect 35437 3587 35495 3593
rect 35437 3553 35449 3587
rect 35483 3584 35495 3587
rect 35866 3584 35894 3624
rect 37918 3612 37924 3624
rect 37976 3612 37982 3664
rect 36814 3584 36820 3596
rect 35483 3556 35894 3584
rect 36775 3556 36820 3584
rect 35483 3553 35495 3556
rect 35437 3547 35495 3553
rect 36814 3544 36820 3556
rect 36872 3544 36878 3596
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 23201 3519 23259 3525
rect 22612 3488 22657 3516
rect 22612 3476 22618 3488
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 23382 3516 23388 3528
rect 23247 3488 23388 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 24670 3516 24676 3528
rect 24631 3488 24676 3516
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 30561 3519 30619 3525
rect 30561 3485 30573 3519
rect 30607 3516 30619 3519
rect 31021 3519 31079 3525
rect 31021 3516 31033 3519
rect 30607 3488 31033 3516
rect 30607 3485 30619 3488
rect 30561 3479 30619 3485
rect 31021 3485 31033 3488
rect 31067 3485 31079 3519
rect 31021 3479 31079 3485
rect 33505 3519 33563 3525
rect 33505 3485 33517 3519
rect 33551 3516 33563 3519
rect 33594 3516 33600 3528
rect 33551 3488 33600 3516
rect 33551 3485 33563 3488
rect 33505 3479 33563 3485
rect 8864 3420 17632 3448
rect 24302 3408 24308 3460
rect 24360 3448 24366 3460
rect 24360 3420 24900 3448
rect 24360 3408 24366 3420
rect 5132 3352 6914 3380
rect 7653 3383 7711 3389
rect 5132 3340 5138 3352
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 9122 3380 9128 3392
rect 7699 3352 9128 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 14458 3340 14464 3392
rect 14516 3380 14522 3392
rect 14553 3383 14611 3389
rect 14553 3380 14565 3383
rect 14516 3352 14565 3380
rect 14516 3340 14522 3352
rect 14553 3349 14565 3352
rect 14599 3349 14611 3383
rect 14553 3343 14611 3349
rect 16393 3383 16451 3389
rect 16393 3349 16405 3383
rect 16439 3380 16451 3383
rect 16850 3380 16856 3392
rect 16439 3352 16856 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 16850 3340 16856 3352
rect 16908 3340 16914 3392
rect 17681 3383 17739 3389
rect 17681 3349 17693 3383
rect 17727 3380 17739 3383
rect 19150 3380 19156 3392
rect 17727 3352 19156 3380
rect 17727 3349 17739 3352
rect 17681 3343 17739 3349
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 19484 3352 19625 3380
rect 19484 3340 19490 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 24762 3380 24768 3392
rect 24723 3352 24768 3380
rect 19613 3343 19671 3349
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 24872 3380 24900 3420
rect 30742 3408 30748 3460
rect 30800 3448 30806 3460
rect 33520 3448 33548 3479
rect 33594 3476 33600 3488
rect 33652 3476 33658 3528
rect 33965 3519 34023 3525
rect 33965 3485 33977 3519
rect 34011 3516 34023 3519
rect 34698 3516 34704 3528
rect 34011 3488 34704 3516
rect 34011 3485 34023 3488
rect 33965 3479 34023 3485
rect 30800 3420 33548 3448
rect 30800 3408 30806 3420
rect 33980 3380 34008 3479
rect 34698 3476 34704 3488
rect 34756 3476 34762 3528
rect 34793 3519 34851 3525
rect 34793 3485 34805 3519
rect 34839 3485 34851 3519
rect 37734 3516 37740 3528
rect 37695 3488 37740 3516
rect 34793 3479 34851 3485
rect 34422 3408 34428 3460
rect 34480 3448 34486 3460
rect 34808 3448 34836 3479
rect 37734 3476 37740 3488
rect 37792 3476 37798 3528
rect 34480 3420 34836 3448
rect 34885 3451 34943 3457
rect 34480 3408 34486 3420
rect 34885 3417 34897 3451
rect 34931 3448 34943 3451
rect 35621 3451 35679 3457
rect 35621 3448 35633 3451
rect 34931 3420 35633 3448
rect 34931 3417 34943 3420
rect 34885 3411 34943 3417
rect 35621 3417 35633 3420
rect 35667 3417 35679 3451
rect 35621 3411 35679 3417
rect 37366 3408 37372 3460
rect 37424 3448 37430 3460
rect 38194 3448 38200 3460
rect 37424 3420 38200 3448
rect 37424 3408 37430 3420
rect 38194 3408 38200 3420
rect 38252 3408 38258 3460
rect 24872 3352 34008 3380
rect 34057 3383 34115 3389
rect 34057 3349 34069 3383
rect 34103 3380 34115 3383
rect 35066 3380 35072 3392
rect 34103 3352 35072 3380
rect 34103 3349 34115 3352
rect 34057 3343 34115 3349
rect 35066 3340 35072 3352
rect 35124 3340 35130 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 4338 3176 4344 3188
rect 4299 3148 4344 3176
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 16298 3176 16304 3188
rect 5684 3148 16304 3176
rect 5684 3136 5690 3148
rect 16298 3136 16304 3148
rect 16356 3176 16362 3188
rect 30837 3179 30895 3185
rect 16356 3148 24440 3176
rect 16356 3136 16362 3148
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 5721 3111 5779 3117
rect 5721 3077 5733 3111
rect 5767 3108 5779 3111
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 5767 3080 6561 3108
rect 5767 3077 5779 3080
rect 5721 3071 5779 3077
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 9214 3108 9220 3120
rect 9175 3080 9220 3108
rect 6549 3071 6607 3077
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 14458 3108 14464 3120
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 16850 3108 16856 3120
rect 16811 3080 16856 3108
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 19150 3108 19156 3120
rect 19111 3080 19156 3108
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 24302 3108 24308 3120
rect 20364 3080 24308 3108
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4212 3012 4445 3040
rect 4212 3000 4218 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 5074 3040 5080 3052
rect 5035 3012 5080 3040
rect 4433 3003 4491 3009
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 4448 2972 4476 3003
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5626 3040 5632 3052
rect 5587 3012 5632 3040
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 9030 3040 9036 3052
rect 8991 3012 9036 3040
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14274 3040 14280 3052
rect 13872 3012 13917 3040
rect 14235 3012 14280 3040
rect 13872 3000 13878 3012
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 18966 3040 18972 3052
rect 18927 3012 18972 3040
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 4614 2972 4620 2984
rect 4448 2944 4620 2972
rect 4614 2932 4620 2944
rect 4672 2972 4678 2984
rect 4672 2944 6500 2972
rect 4672 2932 4678 2944
rect 3878 2864 3884 2916
rect 3936 2904 3942 2916
rect 6472 2904 6500 2944
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6696 2944 6837 2972
rect 6696 2932 6702 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 9674 2972 9680 2984
rect 9635 2944 9680 2972
rect 6825 2935 6883 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 13357 2975 13415 2981
rect 13357 2941 13369 2975
rect 13403 2941 13415 2975
rect 13630 2972 13636 2984
rect 13591 2944 13636 2972
rect 13357 2935 13415 2941
rect 13372 2904 13400 2935
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 14826 2972 14832 2984
rect 14787 2944 14832 2972
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 16666 2972 16672 2984
rect 16627 2944 16672 2972
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 16776 2944 17141 2972
rect 16776 2916 16804 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 18046 2932 18052 2984
rect 18104 2972 18110 2984
rect 19429 2975 19487 2981
rect 19429 2972 19441 2975
rect 18104 2944 19441 2972
rect 18104 2932 18110 2944
rect 19429 2941 19441 2944
rect 19475 2941 19487 2975
rect 19429 2935 19487 2941
rect 13538 2904 13544 2916
rect 3936 2876 6408 2904
rect 6472 2876 11744 2904
rect 13372 2876 13544 2904
rect 3936 2864 3942 2876
rect 4985 2839 5043 2845
rect 4985 2805 4997 2839
rect 5031 2836 5043 2839
rect 5442 2836 5448 2848
rect 5031 2808 5448 2836
rect 5031 2805 5043 2808
rect 4985 2799 5043 2805
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 6380 2836 6408 2876
rect 6822 2836 6828 2848
rect 6380 2808 6828 2836
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 11716 2836 11744 2876
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 16758 2864 16764 2916
rect 16816 2864 16822 2916
rect 20364 2836 20392 3080
rect 24302 3068 24308 3080
rect 24360 3068 24366 3120
rect 21821 2975 21879 2981
rect 21821 2941 21833 2975
rect 21867 2941 21879 2975
rect 22002 2972 22008 2984
rect 21963 2944 22008 2972
rect 21821 2935 21879 2941
rect 21836 2904 21864 2935
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 22557 2975 22615 2981
rect 22557 2941 22569 2975
rect 22603 2941 22615 2975
rect 22557 2935 22615 2941
rect 22462 2904 22468 2916
rect 21836 2876 22468 2904
rect 22462 2864 22468 2876
rect 22520 2864 22526 2916
rect 11716 2808 20392 2836
rect 21910 2796 21916 2848
rect 21968 2836 21974 2848
rect 22572 2836 22600 2935
rect 24412 2904 24440 3148
rect 30837 3145 30849 3179
rect 30883 3176 30895 3179
rect 32398 3176 32404 3188
rect 30883 3148 32404 3176
rect 30883 3145 30895 3148
rect 30837 3139 30895 3145
rect 32398 3136 32404 3148
rect 32456 3136 32462 3188
rect 32490 3136 32496 3188
rect 32548 3176 32554 3188
rect 32548 3148 37412 3176
rect 32548 3136 32554 3148
rect 24762 3108 24768 3120
rect 24723 3080 24768 3108
rect 24762 3068 24768 3080
rect 24820 3068 24826 3120
rect 31481 3111 31539 3117
rect 31481 3077 31493 3111
rect 31527 3108 31539 3111
rect 32309 3111 32367 3117
rect 32309 3108 32321 3111
rect 31527 3080 32321 3108
rect 31527 3077 31539 3080
rect 31481 3071 31539 3077
rect 32309 3077 32321 3080
rect 32355 3077 32367 3111
rect 35066 3108 35072 3120
rect 35027 3080 35072 3108
rect 32309 3071 32367 3077
rect 35066 3068 35072 3080
rect 35124 3068 35130 3120
rect 30742 3040 30748 3052
rect 30703 3012 30748 3040
rect 30742 3000 30748 3012
rect 30800 3000 30806 3052
rect 31386 3040 31392 3052
rect 31347 3012 31392 3040
rect 31386 3000 31392 3012
rect 31444 3000 31450 3052
rect 34790 3000 34796 3052
rect 34848 3040 34854 3052
rect 37384 3049 37412 3148
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 34848 3012 34897 3040
rect 34848 3000 34854 3012
rect 34885 3009 34897 3012
rect 34931 3009 34943 3043
rect 34885 3003 34943 3009
rect 37369 3043 37427 3049
rect 37369 3009 37381 3043
rect 37415 3040 37427 3043
rect 37458 3040 37464 3052
rect 37415 3012 37464 3040
rect 37415 3009 37427 3012
rect 37369 3003 37427 3009
rect 37458 3000 37464 3012
rect 37516 3000 37522 3052
rect 24578 2972 24584 2984
rect 24539 2944 24584 2972
rect 24578 2932 24584 2944
rect 24636 2932 24642 2984
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 32122 2972 32128 2984
rect 32083 2944 32128 2972
rect 32122 2932 32128 2944
rect 32180 2932 32186 2984
rect 32585 2975 32643 2981
rect 32585 2972 32597 2975
rect 32232 2944 32597 2972
rect 32232 2916 32260 2944
rect 32585 2941 32597 2944
rect 32631 2941 32643 2975
rect 35434 2972 35440 2984
rect 35395 2944 35440 2972
rect 32585 2935 32643 2941
rect 35434 2932 35440 2944
rect 35492 2932 35498 2984
rect 24412 2876 31754 2904
rect 21968 2808 22600 2836
rect 31726 2836 31754 2876
rect 32214 2864 32220 2916
rect 32272 2864 32278 2916
rect 34422 2836 34428 2848
rect 31726 2808 34428 2836
rect 21968 2796 21974 2808
rect 34422 2796 34428 2808
rect 34480 2796 34486 2848
rect 36538 2796 36544 2848
rect 36596 2836 36602 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36596 2808 37473 2836
rect 36596 2796 36602 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 13630 2632 13636 2644
rect 13311 2604 13636 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 16666 2632 16672 2644
rect 16627 2604 16672 2632
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 21913 2635 21971 2641
rect 21913 2601 21925 2635
rect 21959 2632 21971 2635
rect 22002 2632 22008 2644
rect 21959 2604 22008 2632
rect 21959 2601 21971 2604
rect 21913 2595 21971 2601
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22462 2632 22468 2644
rect 22423 2604 22468 2632
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 22554 2592 22560 2644
rect 22612 2632 22618 2644
rect 23109 2635 23167 2641
rect 23109 2632 23121 2635
rect 22612 2604 23121 2632
rect 22612 2592 22618 2604
rect 23109 2601 23121 2604
rect 23155 2601 23167 2635
rect 23109 2595 23167 2601
rect 24578 2592 24584 2644
rect 24636 2632 24642 2644
rect 24673 2635 24731 2641
rect 24673 2632 24685 2635
rect 24636 2604 24685 2632
rect 24636 2592 24642 2604
rect 24673 2601 24685 2604
rect 24719 2601 24731 2635
rect 24673 2595 24731 2601
rect 31573 2635 31631 2641
rect 31573 2601 31585 2635
rect 31619 2632 31631 2635
rect 32122 2632 32128 2644
rect 31619 2604 32128 2632
rect 31619 2601 31631 2604
rect 31573 2595 31631 2601
rect 32122 2592 32128 2604
rect 32180 2592 32186 2644
rect 37918 2632 37924 2644
rect 33704 2604 37780 2632
rect 37879 2604 37924 2632
rect 19426 2524 19432 2576
rect 19484 2524 19490 2576
rect 30929 2567 30987 2573
rect 30929 2533 30941 2567
rect 30975 2564 30987 2567
rect 31754 2564 31760 2576
rect 30975 2536 31760 2564
rect 30975 2533 30987 2536
rect 30929 2527 30987 2533
rect 31754 2524 31760 2536
rect 31812 2524 31818 2576
rect 3050 2496 3056 2508
rect 3011 2468 3056 2496
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 4062 2496 4068 2508
rect 3283 2468 4068 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 5442 2496 5448 2508
rect 5403 2468 5448 2496
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 5994 2496 6000 2508
rect 5675 2468 6000 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6270 2456 6276 2508
rect 6328 2496 6334 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 6328 2468 6377 2496
rect 6328 2456 6334 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6365 2459 6423 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6822 2496 6828 2508
rect 6783 2468 6828 2496
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 8386 2456 8392 2508
rect 8444 2496 8450 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 8444 2468 9413 2496
rect 8444 2456 8450 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 19444 2496 19472 2524
rect 19521 2499 19579 2505
rect 19521 2496 19533 2499
rect 19444 2468 19533 2496
rect 9401 2459 9459 2465
rect 19521 2465 19533 2468
rect 19567 2465 19579 2499
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19521 2459 19579 2465
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 33704 2505 33732 2604
rect 37369 2567 37427 2573
rect 37369 2564 37381 2567
rect 36372 2536 37381 2564
rect 33689 2499 33747 2505
rect 33689 2465 33701 2499
rect 33735 2465 33747 2499
rect 33689 2459 33747 2465
rect 33965 2499 34023 2505
rect 33965 2465 33977 2499
rect 34011 2496 34023 2499
rect 36372 2496 36400 2536
rect 37369 2533 37381 2536
rect 37415 2533 37427 2567
rect 37752 2564 37780 2604
rect 37918 2592 37924 2604
rect 37976 2592 37982 2644
rect 38010 2564 38016 2576
rect 37752 2536 38016 2564
rect 37369 2527 37427 2533
rect 38010 2524 38016 2536
rect 38068 2524 38074 2576
rect 36538 2496 36544 2508
rect 34011 2468 36400 2496
rect 36499 2468 36544 2496
rect 34011 2465 34023 2468
rect 33965 2459 34023 2465
rect 36538 2456 36544 2468
rect 36596 2456 36602 2508
rect 36722 2496 36728 2508
rect 36683 2468 36728 2496
rect 36722 2456 36728 2468
rect 36780 2456 36786 2508
rect 8938 2428 8944 2440
rect 8899 2400 8944 2428
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 13354 2388 13360 2400
rect 13412 2428 13418 2440
rect 18693 2431 18751 2437
rect 13412 2400 16574 2428
rect 13412 2388 13418 2400
rect 1394 2360 1400 2372
rect 1355 2332 1400 2360
rect 1394 2320 1400 2332
rect 1452 2320 1458 2372
rect 3789 2363 3847 2369
rect 3789 2360 3801 2363
rect 3252 2332 3801 2360
rect 3252 2304 3280 2332
rect 3789 2329 3801 2332
rect 3835 2329 3847 2363
rect 9122 2360 9128 2372
rect 9083 2332 9128 2360
rect 3789 2323 3847 2329
rect 9122 2320 9128 2332
rect 9180 2320 9186 2372
rect 16546 2360 16574 2400
rect 18693 2397 18705 2431
rect 18739 2428 18751 2431
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 18739 2400 19349 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 19337 2391 19395 2397
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34514 2428 34520 2440
rect 34195 2400 34520 2428
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 21542 2360 21548 2372
rect 16546 2332 21548 2360
rect 21542 2320 21548 2332
rect 21600 2360 21606 2372
rect 21836 2360 21864 2391
rect 34514 2388 34520 2400
rect 34572 2388 34578 2440
rect 36906 2388 36912 2440
rect 36964 2428 36970 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36964 2400 37289 2428
rect 36964 2388 36970 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 21600 2332 21864 2360
rect 34885 2363 34943 2369
rect 21600 2320 21606 2332
rect 34885 2329 34897 2363
rect 34931 2360 34943 2363
rect 35158 2360 35164 2372
rect 34931 2332 35164 2360
rect 34931 2329 34943 2332
rect 34885 2323 34943 2329
rect 35158 2320 35164 2332
rect 35216 2320 35222 2372
rect 3234 2252 3240 2304
rect 3292 2252 3298 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 11520 37340 11572 37392
rect 34888 37340 34940 37392
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 2136 37204 2188 37256
rect 1952 37136 2004 37188
rect 2044 37068 2096 37120
rect 2228 37111 2280 37120
rect 2228 37077 2237 37111
rect 2237 37077 2271 37111
rect 2271 37077 2280 37111
rect 2228 37068 2280 37077
rect 3056 37068 3108 37120
rect 5632 37247 5684 37256
rect 5632 37213 5641 37247
rect 5641 37213 5675 37247
rect 5675 37213 5684 37247
rect 6644 37247 6696 37256
rect 5632 37204 5684 37213
rect 6644 37213 6653 37247
rect 6653 37213 6687 37247
rect 6687 37213 6696 37247
rect 6644 37204 6696 37213
rect 7748 37247 7800 37256
rect 7748 37213 7757 37247
rect 7757 37213 7791 37247
rect 7791 37213 7800 37247
rect 7748 37204 7800 37213
rect 9772 37247 9824 37256
rect 9772 37213 9781 37247
rect 9781 37213 9815 37247
rect 9815 37213 9824 37247
rect 9772 37204 9824 37213
rect 11704 37272 11756 37324
rect 16120 37272 16172 37324
rect 20628 37315 20680 37324
rect 17684 37247 17736 37256
rect 10876 37136 10928 37188
rect 12164 37136 12216 37188
rect 17684 37213 17693 37247
rect 17693 37213 17727 37247
rect 17727 37213 17736 37247
rect 17684 37204 17736 37213
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 20628 37281 20637 37315
rect 20637 37281 20671 37315
rect 20671 37281 20680 37315
rect 20628 37272 20680 37281
rect 27252 37315 27304 37324
rect 27252 37281 27261 37315
rect 27261 37281 27295 37315
rect 27295 37281 27304 37315
rect 27252 37272 27304 37281
rect 21824 37247 21876 37256
rect 21824 37213 21833 37247
rect 21833 37213 21867 37247
rect 21867 37213 21876 37247
rect 21824 37204 21876 37213
rect 23112 37204 23164 37256
rect 23664 37247 23716 37256
rect 23664 37213 23673 37247
rect 23673 37213 23707 37247
rect 23707 37213 23716 37247
rect 23664 37204 23716 37213
rect 24124 37204 24176 37256
rect 25412 37247 25464 37256
rect 25412 37213 25421 37247
rect 25421 37213 25455 37247
rect 25455 37213 25464 37247
rect 25412 37204 25464 37213
rect 25780 37204 25832 37256
rect 26148 37204 26200 37256
rect 36728 37315 36780 37324
rect 36728 37281 36737 37315
rect 36737 37281 36771 37315
rect 36771 37281 36780 37315
rect 36728 37272 36780 37281
rect 37280 37247 37332 37256
rect 37280 37213 37289 37247
rect 37289 37213 37323 37247
rect 37323 37213 37332 37247
rect 37280 37204 37332 37213
rect 37924 37247 37976 37256
rect 37924 37213 37933 37247
rect 37933 37213 37967 37247
rect 37967 37213 37976 37247
rect 37924 37204 37976 37213
rect 5816 37068 5868 37120
rect 6460 37111 6512 37120
rect 6460 37077 6469 37111
rect 6469 37077 6503 37111
rect 6503 37077 6512 37111
rect 6460 37068 6512 37077
rect 7288 37068 7340 37120
rect 12716 37068 12768 37120
rect 14188 37111 14240 37120
rect 14188 37077 14197 37111
rect 14197 37077 14231 37111
rect 14231 37077 14240 37111
rect 14188 37068 14240 37077
rect 20076 37136 20128 37188
rect 22376 37136 22428 37188
rect 29552 37136 29604 37188
rect 29644 37136 29696 37188
rect 30932 37136 30984 37188
rect 34796 37136 34848 37188
rect 36544 37136 36596 37188
rect 21732 37068 21784 37120
rect 21916 37111 21968 37120
rect 21916 37077 21925 37111
rect 21925 37077 21959 37111
rect 21959 37077 21968 37111
rect 21916 37068 21968 37077
rect 22836 37068 22888 37120
rect 25964 37111 26016 37120
rect 25964 37077 25973 37111
rect 25973 37077 26007 37111
rect 26007 37077 26016 37111
rect 25964 37068 26016 37077
rect 28724 37111 28776 37120
rect 28724 37077 28733 37111
rect 28733 37077 28767 37111
rect 28767 37077 28776 37111
rect 28724 37068 28776 37077
rect 35900 37068 35952 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2044 36864 2096 36916
rect 5724 36864 5776 36916
rect 6644 36864 6696 36916
rect 10876 36907 10928 36916
rect 10876 36873 10885 36907
rect 10885 36873 10919 36907
rect 10919 36873 10928 36907
rect 10876 36864 10928 36873
rect 1584 36839 1636 36848
rect 1584 36805 1593 36839
rect 1593 36805 1627 36839
rect 1627 36805 1636 36839
rect 1584 36796 1636 36805
rect 2228 36796 2280 36848
rect 3884 36839 3936 36848
rect 3884 36805 3893 36839
rect 3893 36805 3927 36839
rect 3927 36805 3936 36839
rect 3884 36796 3936 36805
rect 7748 36796 7800 36848
rect 10508 36796 10560 36848
rect 12624 36864 12676 36916
rect 12716 36864 12768 36916
rect 23112 36864 23164 36916
rect 25780 36864 25832 36916
rect 6460 36771 6512 36780
rect 6460 36737 6469 36771
rect 6469 36737 6503 36771
rect 6503 36737 6512 36771
rect 6460 36728 6512 36737
rect 7196 36771 7248 36780
rect 7196 36737 7205 36771
rect 7205 36737 7239 36771
rect 7239 36737 7248 36771
rect 7196 36728 7248 36737
rect 10416 36728 10468 36780
rect 12072 36796 12124 36848
rect 12256 36796 12308 36848
rect 11520 36771 11572 36780
rect 11520 36737 11529 36771
rect 11529 36737 11563 36771
rect 11563 36737 11572 36771
rect 11520 36728 11572 36737
rect 3424 36703 3476 36712
rect 3424 36669 3433 36703
rect 3433 36669 3467 36703
rect 3467 36669 3476 36703
rect 3424 36660 3476 36669
rect 5540 36703 5592 36712
rect 5540 36669 5549 36703
rect 5549 36669 5583 36703
rect 5583 36669 5592 36703
rect 5540 36660 5592 36669
rect 8392 36703 8444 36712
rect 8392 36669 8401 36703
rect 8401 36669 8435 36703
rect 8435 36669 8444 36703
rect 8392 36660 8444 36669
rect 9036 36660 9088 36712
rect 11704 36703 11756 36712
rect 11704 36669 11713 36703
rect 11713 36669 11747 36703
rect 11747 36669 11756 36703
rect 11704 36660 11756 36669
rect 9680 36592 9732 36644
rect 10968 36592 11020 36644
rect 12072 36660 12124 36712
rect 16120 36771 16172 36780
rect 16120 36737 16129 36771
rect 16129 36737 16163 36771
rect 16163 36737 16172 36771
rect 17132 36771 17184 36780
rect 16120 36728 16172 36737
rect 17132 36737 17141 36771
rect 17141 36737 17175 36771
rect 17175 36737 17184 36771
rect 17132 36728 17184 36737
rect 17684 36771 17736 36780
rect 17684 36737 17693 36771
rect 17693 36737 17727 36771
rect 17727 36737 17736 36771
rect 17684 36728 17736 36737
rect 17040 36660 17092 36712
rect 17868 36703 17920 36712
rect 17868 36669 17877 36703
rect 17877 36669 17911 36703
rect 17911 36669 17920 36703
rect 17868 36660 17920 36669
rect 18052 36660 18104 36712
rect 21272 36796 21324 36848
rect 21180 36771 21232 36780
rect 21180 36737 21189 36771
rect 21189 36737 21223 36771
rect 21223 36737 21232 36771
rect 21180 36728 21232 36737
rect 23664 36771 23716 36780
rect 23664 36737 23673 36771
rect 23673 36737 23707 36771
rect 23707 36737 23716 36771
rect 24124 36771 24176 36780
rect 23664 36728 23716 36737
rect 24124 36737 24133 36771
rect 24133 36737 24167 36771
rect 24167 36737 24176 36771
rect 24124 36728 24176 36737
rect 28264 36728 28316 36780
rect 34888 36771 34940 36780
rect 21916 36660 21968 36712
rect 24492 36660 24544 36712
rect 24584 36703 24636 36712
rect 24584 36669 24593 36703
rect 24593 36669 24627 36703
rect 24627 36669 24636 36703
rect 34888 36737 34897 36771
rect 34897 36737 34931 36771
rect 34931 36737 34940 36771
rect 34888 36728 34940 36737
rect 37188 36728 37240 36780
rect 38568 36728 38620 36780
rect 24584 36660 24636 36669
rect 10692 36524 10744 36576
rect 26792 36592 26844 36644
rect 16948 36524 17000 36576
rect 17132 36524 17184 36576
rect 19432 36524 19484 36576
rect 21640 36524 21692 36576
rect 29000 36660 29052 36712
rect 30196 36660 30248 36712
rect 32404 36703 32456 36712
rect 29736 36592 29788 36644
rect 32404 36669 32413 36703
rect 32413 36669 32447 36703
rect 32447 36669 32456 36703
rect 32404 36660 32456 36669
rect 32588 36703 32640 36712
rect 32588 36669 32597 36703
rect 32597 36669 32631 36703
rect 32631 36669 32640 36703
rect 32588 36660 32640 36669
rect 32864 36703 32916 36712
rect 32864 36669 32873 36703
rect 32873 36669 32907 36703
rect 32907 36669 32916 36703
rect 32864 36660 32916 36669
rect 27804 36524 27856 36576
rect 27988 36524 28040 36576
rect 31668 36524 31720 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 9036 36363 9088 36372
rect 9036 36329 9045 36363
rect 9045 36329 9079 36363
rect 9079 36329 9088 36363
rect 9036 36320 9088 36329
rect 9864 36320 9916 36372
rect 10416 36320 10468 36372
rect 12624 36320 12676 36372
rect 17040 36363 17092 36372
rect 2136 36252 2188 36304
rect 17040 36329 17049 36363
rect 17049 36329 17083 36363
rect 17083 36329 17092 36363
rect 17040 36320 17092 36329
rect 17868 36363 17920 36372
rect 17868 36329 17877 36363
rect 17877 36329 17911 36363
rect 17911 36329 17920 36363
rect 17868 36320 17920 36329
rect 20076 36320 20128 36372
rect 24492 36363 24544 36372
rect 24492 36329 24501 36363
rect 24501 36329 24535 36363
rect 24535 36329 24544 36363
rect 24492 36320 24544 36329
rect 29644 36363 29696 36372
rect 29644 36329 29653 36363
rect 29653 36329 29687 36363
rect 29687 36329 29696 36363
rect 29644 36320 29696 36329
rect 30196 36363 30248 36372
rect 30196 36329 30205 36363
rect 30205 36329 30239 36363
rect 30239 36329 30248 36363
rect 30196 36320 30248 36329
rect 34796 36363 34848 36372
rect 34796 36329 34805 36363
rect 34805 36329 34839 36363
rect 34839 36329 34848 36363
rect 34796 36320 34848 36329
rect 1308 36184 1360 36236
rect 3056 36227 3108 36236
rect 3056 36193 3065 36227
rect 3065 36193 3099 36227
rect 3099 36193 3108 36227
rect 3056 36184 3108 36193
rect 4620 36227 4672 36236
rect 4620 36193 4629 36227
rect 4629 36193 4663 36227
rect 4663 36193 4672 36227
rect 4620 36184 4672 36193
rect 9772 36227 9824 36236
rect 9772 36193 9781 36227
rect 9781 36193 9815 36227
rect 9815 36193 9824 36227
rect 9772 36184 9824 36193
rect 10324 36227 10376 36236
rect 10324 36193 10333 36227
rect 10333 36193 10367 36227
rect 10367 36193 10376 36227
rect 10324 36184 10376 36193
rect 18512 36252 18564 36304
rect 22008 36252 22060 36304
rect 16304 36184 16356 36236
rect 18696 36184 18748 36236
rect 19984 36227 20036 36236
rect 19984 36193 19993 36227
rect 19993 36193 20027 36227
rect 20027 36193 20036 36227
rect 19984 36184 20036 36193
rect 25412 36184 25464 36236
rect 25964 36227 26016 36236
rect 25964 36193 25973 36227
rect 25973 36193 26007 36227
rect 26007 36193 26016 36227
rect 25964 36184 26016 36193
rect 26424 36227 26476 36236
rect 26424 36193 26433 36227
rect 26433 36193 26467 36227
rect 26467 36193 26476 36227
rect 26424 36184 26476 36193
rect 31668 36227 31720 36236
rect 31668 36193 31677 36227
rect 31677 36193 31711 36227
rect 31711 36193 31720 36227
rect 31668 36184 31720 36193
rect 32220 36227 32272 36236
rect 32220 36193 32229 36227
rect 32229 36193 32263 36227
rect 32263 36193 32272 36227
rect 32220 36184 32272 36193
rect 38108 36227 38160 36236
rect 38108 36193 38117 36227
rect 38117 36193 38151 36227
rect 38151 36193 38160 36227
rect 38108 36184 38160 36193
rect 6460 36159 6512 36168
rect 2964 36048 3016 36100
rect 6460 36125 6469 36159
rect 6469 36125 6503 36159
rect 6503 36125 6512 36159
rect 6460 36116 6512 36125
rect 8852 36116 8904 36168
rect 12164 36159 12216 36168
rect 12164 36125 12173 36159
rect 12173 36125 12207 36159
rect 12207 36125 12216 36159
rect 12164 36116 12216 36125
rect 13544 36116 13596 36168
rect 16396 36116 16448 36168
rect 16488 36159 16540 36168
rect 16488 36125 16497 36159
rect 16497 36125 16531 36159
rect 16531 36125 16540 36159
rect 16488 36116 16540 36125
rect 17776 36159 17828 36168
rect 4620 36048 4672 36100
rect 5816 36048 5868 36100
rect 9772 36048 9824 36100
rect 9956 36091 10008 36100
rect 9956 36057 9965 36091
rect 9965 36057 9999 36091
rect 9999 36057 10008 36091
rect 9956 36048 10008 36057
rect 12532 36048 12584 36100
rect 13360 36048 13412 36100
rect 14188 36048 14240 36100
rect 15568 36091 15620 36100
rect 15568 36057 15577 36091
rect 15577 36057 15611 36091
rect 15611 36057 15620 36091
rect 15568 36048 15620 36057
rect 9864 35980 9916 36032
rect 10692 35980 10744 36032
rect 12440 35980 12492 36032
rect 14096 36023 14148 36032
rect 14096 35989 14105 36023
rect 14105 35989 14139 36023
rect 14139 35989 14148 36023
rect 14096 35980 14148 35989
rect 15660 35980 15712 36032
rect 17776 36125 17785 36159
rect 17785 36125 17819 36159
rect 17819 36125 17828 36159
rect 17776 36116 17828 36125
rect 18512 36159 18564 36168
rect 18512 36125 18521 36159
rect 18521 36125 18555 36159
rect 18555 36125 18564 36159
rect 18512 36116 18564 36125
rect 21180 36116 21232 36168
rect 22652 36116 22704 36168
rect 24584 36159 24636 36168
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 25320 36116 25372 36168
rect 22376 36091 22428 36100
rect 22376 36057 22385 36091
rect 22385 36057 22419 36091
rect 22419 36057 22428 36091
rect 22376 36048 22428 36057
rect 28540 36116 28592 36168
rect 29000 36116 29052 36168
rect 34612 36116 34664 36168
rect 34704 36159 34756 36168
rect 34704 36125 34713 36159
rect 34713 36125 34747 36159
rect 34747 36125 34756 36159
rect 34704 36116 34756 36125
rect 28816 36048 28868 36100
rect 31852 36091 31904 36100
rect 31852 36057 31861 36091
rect 31861 36057 31895 36091
rect 31895 36057 31904 36091
rect 31852 36048 31904 36057
rect 37464 36048 37516 36100
rect 20904 35980 20956 36032
rect 25044 35980 25096 36032
rect 28448 35980 28500 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 5540 35776 5592 35828
rect 9128 35776 9180 35828
rect 9680 35776 9732 35828
rect 9956 35776 10008 35828
rect 11704 35776 11756 35828
rect 15568 35776 15620 35828
rect 21732 35776 21784 35828
rect 27252 35776 27304 35828
rect 29552 35776 29604 35828
rect 31852 35776 31904 35828
rect 32588 35776 32640 35828
rect 37464 35819 37516 35828
rect 37464 35785 37473 35819
rect 37473 35785 37507 35819
rect 37507 35785 37516 35819
rect 37464 35776 37516 35785
rect 7288 35708 7340 35760
rect 12532 35708 12584 35760
rect 21364 35708 21416 35760
rect 35900 35708 35952 35760
rect 38016 35708 38068 35760
rect 6460 35683 6512 35692
rect 1768 35615 1820 35624
rect 1768 35581 1777 35615
rect 1777 35581 1811 35615
rect 1811 35581 1820 35615
rect 1768 35572 1820 35581
rect 2228 35572 2280 35624
rect 2780 35615 2832 35624
rect 2780 35581 2789 35615
rect 2789 35581 2823 35615
rect 2823 35581 2832 35615
rect 2780 35572 2832 35581
rect 6460 35649 6469 35683
rect 6469 35649 6503 35683
rect 6503 35649 6512 35683
rect 6460 35640 6512 35649
rect 8392 35683 8444 35692
rect 8392 35649 8401 35683
rect 8401 35649 8435 35683
rect 8435 35649 8444 35683
rect 8392 35640 8444 35649
rect 9864 35640 9916 35692
rect 10508 35683 10560 35692
rect 10508 35649 10517 35683
rect 10517 35649 10551 35683
rect 10551 35649 10560 35683
rect 10508 35640 10560 35649
rect 14096 35640 14148 35692
rect 14372 35683 14424 35692
rect 14372 35649 14389 35683
rect 14389 35649 14424 35683
rect 14372 35640 14424 35649
rect 14464 35683 14516 35692
rect 14464 35649 14473 35683
rect 14473 35649 14507 35683
rect 14507 35649 14516 35683
rect 14464 35640 14516 35649
rect 15108 35640 15160 35692
rect 15292 35683 15344 35692
rect 15292 35649 15301 35683
rect 15301 35649 15335 35683
rect 15335 35649 15344 35683
rect 15292 35640 15344 35649
rect 15936 35683 15988 35692
rect 6000 35572 6052 35624
rect 7196 35615 7248 35624
rect 7196 35581 7205 35615
rect 7205 35581 7239 35615
rect 7239 35581 7248 35615
rect 7196 35572 7248 35581
rect 11520 35572 11572 35624
rect 11980 35615 12032 35624
rect 11980 35581 11989 35615
rect 11989 35581 12023 35615
rect 12023 35581 12032 35615
rect 11980 35572 12032 35581
rect 13820 35572 13872 35624
rect 15936 35649 15945 35683
rect 15945 35649 15979 35683
rect 15979 35649 15988 35683
rect 15936 35640 15988 35649
rect 16396 35640 16448 35692
rect 19340 35640 19392 35692
rect 19524 35683 19576 35692
rect 19524 35649 19533 35683
rect 19533 35649 19567 35683
rect 19567 35649 19576 35683
rect 19524 35640 19576 35649
rect 20260 35640 20312 35692
rect 17684 35572 17736 35624
rect 11244 35436 11296 35488
rect 20720 35640 20772 35692
rect 21180 35640 21232 35692
rect 22008 35683 22060 35692
rect 22008 35649 22017 35683
rect 22017 35649 22051 35683
rect 22051 35649 22060 35683
rect 22008 35640 22060 35649
rect 22652 35683 22704 35692
rect 22652 35649 22661 35683
rect 22661 35649 22695 35683
rect 22695 35649 22704 35683
rect 22652 35640 22704 35649
rect 25504 35640 25556 35692
rect 26976 35640 27028 35692
rect 27344 35683 27396 35692
rect 27344 35649 27353 35683
rect 27353 35649 27387 35683
rect 27387 35649 27396 35683
rect 27344 35640 27396 35649
rect 27804 35683 27856 35692
rect 27804 35649 27813 35683
rect 27813 35649 27847 35683
rect 27847 35649 27856 35683
rect 27804 35640 27856 35649
rect 30104 35683 30156 35692
rect 30104 35649 30113 35683
rect 30113 35649 30147 35683
rect 30147 35649 30156 35683
rect 30104 35640 30156 35649
rect 32220 35640 32272 35692
rect 32588 35640 32640 35692
rect 34612 35640 34664 35692
rect 20812 35615 20864 35624
rect 20812 35581 20821 35615
rect 20821 35581 20855 35615
rect 20855 35581 20864 35615
rect 20812 35572 20864 35581
rect 22836 35615 22888 35624
rect 22836 35581 22845 35615
rect 22845 35581 22879 35615
rect 22879 35581 22888 35615
rect 22836 35572 22888 35581
rect 23204 35615 23256 35624
rect 23204 35581 23213 35615
rect 23213 35581 23247 35615
rect 23247 35581 23256 35615
rect 23204 35572 23256 35581
rect 27988 35615 28040 35624
rect 27988 35581 27997 35615
rect 27997 35581 28031 35615
rect 28031 35581 28040 35615
rect 27988 35572 28040 35581
rect 28356 35615 28408 35624
rect 28356 35581 28365 35615
rect 28365 35581 28399 35615
rect 28399 35581 28408 35615
rect 28356 35572 28408 35581
rect 20996 35504 21048 35556
rect 21824 35504 21876 35556
rect 38384 35640 38436 35692
rect 13544 35436 13596 35488
rect 13636 35436 13688 35488
rect 14372 35436 14424 35488
rect 17040 35436 17092 35488
rect 18328 35436 18380 35488
rect 25136 35479 25188 35488
rect 25136 35445 25145 35479
rect 25145 35445 25179 35479
rect 25179 35445 25188 35479
rect 25136 35436 25188 35445
rect 26240 35436 26292 35488
rect 26884 35436 26936 35488
rect 36728 35436 36780 35488
rect 36820 35436 36872 35488
rect 38016 35436 38068 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4620 35232 4672 35284
rect 11980 35232 12032 35284
rect 12532 35232 12584 35284
rect 15292 35232 15344 35284
rect 17684 35275 17736 35284
rect 17684 35241 17693 35275
rect 17693 35241 17727 35275
rect 17727 35241 17736 35275
rect 17684 35232 17736 35241
rect 19340 35275 19392 35284
rect 19340 35241 19349 35275
rect 19349 35241 19383 35275
rect 19383 35241 19392 35275
rect 19340 35232 19392 35241
rect 24584 35232 24636 35284
rect 27344 35275 27396 35284
rect 2872 35096 2924 35148
rect 10692 35096 10744 35148
rect 3240 35071 3292 35080
rect 3240 35037 3249 35071
rect 3249 35037 3283 35071
rect 3283 35037 3292 35071
rect 3240 35028 3292 35037
rect 5816 35071 5868 35080
rect 5816 35037 5825 35071
rect 5825 35037 5859 35071
rect 5859 35037 5868 35071
rect 5816 35028 5868 35037
rect 6460 35071 6512 35080
rect 6460 35037 6469 35071
rect 6469 35037 6503 35071
rect 6503 35037 6512 35071
rect 6460 35028 6512 35037
rect 8484 35028 8536 35080
rect 11244 35071 11296 35080
rect 11244 35037 11253 35071
rect 11253 35037 11287 35071
rect 11287 35037 11296 35071
rect 11244 35028 11296 35037
rect 12164 35028 12216 35080
rect 12440 35071 12492 35080
rect 12440 35037 12449 35071
rect 12449 35037 12483 35071
rect 12483 35037 12492 35071
rect 12440 35028 12492 35037
rect 2872 34960 2924 35012
rect 5448 35003 5500 35012
rect 5448 34969 5457 35003
rect 5457 34969 5491 35003
rect 5491 34969 5500 35003
rect 5448 34960 5500 34969
rect 6184 34960 6236 35012
rect 8852 34960 8904 35012
rect 10784 34960 10836 35012
rect 11980 34960 12032 35012
rect 12532 35003 12584 35012
rect 12532 34969 12541 35003
rect 12541 34969 12575 35003
rect 12575 34969 12584 35003
rect 12532 34960 12584 34969
rect 14464 35164 14516 35216
rect 16212 35164 16264 35216
rect 14096 35096 14148 35148
rect 13360 35071 13412 35080
rect 13360 35037 13369 35071
rect 13369 35037 13403 35071
rect 13403 35037 13412 35071
rect 13360 35028 13412 35037
rect 13544 35071 13596 35080
rect 13544 35037 13553 35071
rect 13553 35037 13587 35071
rect 13587 35037 13596 35071
rect 13544 35028 13596 35037
rect 13912 35028 13964 35080
rect 10600 34892 10652 34944
rect 10692 34935 10744 34944
rect 10692 34901 10701 34935
rect 10701 34901 10735 34935
rect 10735 34901 10744 34935
rect 11704 34935 11756 34944
rect 10692 34892 10744 34901
rect 11704 34901 11713 34935
rect 11713 34901 11747 34935
rect 11747 34901 11756 34935
rect 11704 34892 11756 34901
rect 11888 34892 11940 34944
rect 12716 34960 12768 35012
rect 14464 34960 14516 35012
rect 15936 35096 15988 35148
rect 15292 35028 15344 35080
rect 16304 35028 16356 35080
rect 18144 35164 18196 35216
rect 18328 35096 18380 35148
rect 24860 35139 24912 35148
rect 24860 35105 24869 35139
rect 24869 35105 24903 35139
rect 24903 35105 24912 35139
rect 24860 35096 24912 35105
rect 26148 35096 26200 35148
rect 19432 35071 19484 35080
rect 15384 35003 15436 35012
rect 15384 34969 15393 35003
rect 15393 34969 15427 35003
rect 15427 34969 15436 35003
rect 19432 35037 19441 35071
rect 19441 35037 19475 35071
rect 19475 35037 19484 35071
rect 19432 35028 19484 35037
rect 20168 35028 20220 35080
rect 20720 35071 20772 35080
rect 20720 35037 20729 35071
rect 20729 35037 20763 35071
rect 20763 35037 20772 35071
rect 20720 35028 20772 35037
rect 15384 34960 15436 34969
rect 17040 34960 17092 35012
rect 13636 34892 13688 34944
rect 13820 34892 13872 34944
rect 15200 34892 15252 34944
rect 15476 34892 15528 34944
rect 16856 34892 16908 34944
rect 17408 35003 17460 35012
rect 17408 34969 17417 35003
rect 17417 34969 17451 35003
rect 17451 34969 17460 35003
rect 18144 35003 18196 35012
rect 17408 34960 17460 34969
rect 18144 34969 18153 35003
rect 18153 34969 18187 35003
rect 18187 34969 18196 35003
rect 18144 34960 18196 34969
rect 18328 35003 18380 35012
rect 18328 34969 18337 35003
rect 18337 34969 18371 35003
rect 18371 34969 18380 35003
rect 18328 34960 18380 34969
rect 21364 35003 21416 35012
rect 21364 34969 21373 35003
rect 21373 34969 21407 35003
rect 21407 34969 21416 35003
rect 21364 34960 21416 34969
rect 23664 34935 23716 34944
rect 23664 34901 23673 34935
rect 23673 34901 23707 34935
rect 23707 34901 23716 34935
rect 23664 34892 23716 34901
rect 26240 35028 26292 35080
rect 25136 35003 25188 35012
rect 25136 34969 25145 35003
rect 25145 34969 25179 35003
rect 25179 34969 25188 35003
rect 25136 34960 25188 34969
rect 25228 34892 25280 34944
rect 26608 34935 26660 34944
rect 26608 34901 26617 34935
rect 26617 34901 26651 34935
rect 26651 34901 26660 34935
rect 26608 34892 26660 34901
rect 27344 35241 27353 35275
rect 27353 35241 27387 35275
rect 27387 35241 27396 35275
rect 27344 35232 27396 35241
rect 28540 35232 28592 35284
rect 32404 35275 32456 35284
rect 32404 35241 32413 35275
rect 32413 35241 32447 35275
rect 32447 35241 32456 35275
rect 32404 35232 32456 35241
rect 36728 35232 36780 35284
rect 37924 35232 37976 35284
rect 27528 35071 27580 35080
rect 27528 35037 27537 35071
rect 27537 35037 27571 35071
rect 27571 35037 27580 35071
rect 27528 35028 27580 35037
rect 28264 35071 28316 35080
rect 28264 35037 28273 35071
rect 28273 35037 28307 35071
rect 28307 35037 28316 35071
rect 28264 35028 28316 35037
rect 28540 35071 28592 35080
rect 28540 35037 28549 35071
rect 28549 35037 28583 35071
rect 28583 35037 28592 35071
rect 28540 35028 28592 35037
rect 37188 35139 37240 35148
rect 37188 35105 37197 35139
rect 37197 35105 37231 35139
rect 37231 35105 37240 35139
rect 37188 35096 37240 35105
rect 29000 35028 29052 35080
rect 29920 35028 29972 35080
rect 31300 35071 31352 35080
rect 31300 35037 31309 35071
rect 31309 35037 31343 35071
rect 31343 35037 31352 35071
rect 31300 35028 31352 35037
rect 36728 35028 36780 35080
rect 38108 35071 38160 35080
rect 38108 35037 38117 35071
rect 38117 35037 38151 35071
rect 38151 35037 38160 35071
rect 38108 35028 38160 35037
rect 28448 35003 28500 35012
rect 28448 34969 28457 35003
rect 28457 34969 28491 35003
rect 28491 34969 28500 35003
rect 28448 34960 28500 34969
rect 37556 34960 37608 35012
rect 31392 34892 31444 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2228 34731 2280 34740
rect 2228 34697 2237 34731
rect 2237 34697 2271 34731
rect 2271 34697 2280 34731
rect 2228 34688 2280 34697
rect 2872 34731 2924 34740
rect 2872 34697 2881 34731
rect 2881 34697 2915 34731
rect 2915 34697 2924 34731
rect 2872 34688 2924 34697
rect 10784 34731 10836 34740
rect 10784 34697 10793 34731
rect 10793 34697 10827 34731
rect 10827 34697 10836 34731
rect 10784 34688 10836 34697
rect 1768 34552 1820 34604
rect 2320 34595 2372 34604
rect 2320 34561 2329 34595
rect 2329 34561 2363 34595
rect 2363 34561 2372 34595
rect 2320 34552 2372 34561
rect 4712 34620 4764 34672
rect 10600 34620 10652 34672
rect 11888 34663 11940 34672
rect 11888 34629 11897 34663
rect 11897 34629 11931 34663
rect 11931 34629 11940 34663
rect 11888 34620 11940 34629
rect 12716 34688 12768 34740
rect 14188 34688 14240 34740
rect 15108 34731 15160 34740
rect 15108 34697 15117 34731
rect 15117 34697 15151 34731
rect 15151 34697 15160 34731
rect 15108 34688 15160 34697
rect 9864 34552 9916 34604
rect 11704 34595 11756 34604
rect 3608 34527 3660 34536
rect 3608 34493 3617 34527
rect 3617 34493 3651 34527
rect 3651 34493 3660 34527
rect 3608 34484 3660 34493
rect 3792 34527 3844 34536
rect 3792 34493 3801 34527
rect 3801 34493 3835 34527
rect 3835 34493 3844 34527
rect 3792 34484 3844 34493
rect 3976 34484 4028 34536
rect 8484 34527 8536 34536
rect 8484 34493 8493 34527
rect 8493 34493 8527 34527
rect 8527 34493 8536 34527
rect 8484 34484 8536 34493
rect 9956 34416 10008 34468
rect 11704 34561 11713 34595
rect 11713 34561 11747 34595
rect 11747 34561 11756 34595
rect 11704 34552 11756 34561
rect 11060 34484 11112 34536
rect 12164 34595 12216 34604
rect 12164 34561 12173 34595
rect 12173 34561 12207 34595
rect 12207 34561 12216 34595
rect 13912 34620 13964 34672
rect 14096 34620 14148 34672
rect 12164 34552 12216 34561
rect 14280 34552 14332 34604
rect 15384 34595 15436 34604
rect 15384 34561 15394 34595
rect 15394 34561 15428 34595
rect 15428 34561 15436 34595
rect 16212 34688 16264 34740
rect 17408 34688 17460 34740
rect 15384 34552 15436 34561
rect 17408 34552 17460 34604
rect 12072 34484 12124 34536
rect 15292 34527 15344 34536
rect 13176 34416 13228 34468
rect 13544 34416 13596 34468
rect 15292 34493 15301 34527
rect 15301 34493 15335 34527
rect 15335 34493 15344 34527
rect 15292 34484 15344 34493
rect 15476 34527 15528 34536
rect 15476 34493 15485 34527
rect 15485 34493 15519 34527
rect 15519 34493 15528 34527
rect 21916 34688 21968 34740
rect 20720 34620 20772 34672
rect 24860 34688 24912 34740
rect 25504 34731 25556 34740
rect 25504 34697 25513 34731
rect 25513 34697 25547 34731
rect 25547 34697 25556 34731
rect 25504 34688 25556 34697
rect 28632 34688 28684 34740
rect 29000 34731 29052 34740
rect 29000 34697 29009 34731
rect 29009 34697 29043 34731
rect 29043 34697 29052 34731
rect 29000 34688 29052 34697
rect 18972 34595 19024 34604
rect 18972 34561 18981 34595
rect 18981 34561 19015 34595
rect 19015 34561 19024 34595
rect 18972 34552 19024 34561
rect 20812 34552 20864 34604
rect 22468 34595 22520 34604
rect 22468 34561 22477 34595
rect 22477 34561 22511 34595
rect 22511 34561 22520 34595
rect 22468 34552 22520 34561
rect 23664 34620 23716 34672
rect 25044 34620 25096 34672
rect 26884 34620 26936 34672
rect 25872 34595 25924 34604
rect 15476 34484 15528 34493
rect 15200 34416 15252 34468
rect 15568 34416 15620 34468
rect 18880 34484 18932 34536
rect 20904 34527 20956 34536
rect 20904 34493 20913 34527
rect 20913 34493 20947 34527
rect 20947 34493 20956 34527
rect 20904 34484 20956 34493
rect 21548 34484 21600 34536
rect 25872 34561 25881 34595
rect 25881 34561 25915 34595
rect 25915 34561 25924 34595
rect 25872 34552 25924 34561
rect 27712 34620 27764 34672
rect 28540 34663 28592 34672
rect 28172 34595 28224 34604
rect 28172 34561 28181 34595
rect 28181 34561 28215 34595
rect 28215 34561 28224 34595
rect 28172 34552 28224 34561
rect 28540 34629 28549 34663
rect 28549 34629 28583 34663
rect 28583 34629 28592 34663
rect 28540 34620 28592 34629
rect 31116 34688 31168 34740
rect 31392 34688 31444 34740
rect 37556 34731 37608 34740
rect 25044 34527 25096 34536
rect 25044 34493 25053 34527
rect 25053 34493 25087 34527
rect 25087 34493 25096 34527
rect 25044 34484 25096 34493
rect 25964 34527 26016 34536
rect 25964 34493 25973 34527
rect 25973 34493 26007 34527
rect 26007 34493 26016 34527
rect 25964 34484 26016 34493
rect 26608 34484 26660 34536
rect 28724 34552 28776 34604
rect 28816 34552 28868 34604
rect 36544 34663 36596 34672
rect 36544 34629 36553 34663
rect 36553 34629 36587 34663
rect 36587 34629 36596 34663
rect 36544 34620 36596 34629
rect 37556 34697 37565 34731
rect 37565 34697 37599 34731
rect 37599 34697 37608 34731
rect 37556 34688 37608 34697
rect 32404 34552 32456 34604
rect 33416 34595 33468 34604
rect 33416 34561 33425 34595
rect 33425 34561 33459 34595
rect 33459 34561 33468 34595
rect 33416 34552 33468 34561
rect 34704 34552 34756 34604
rect 36728 34595 36780 34604
rect 36728 34561 36737 34595
rect 36737 34561 36771 34595
rect 36771 34561 36780 34595
rect 36728 34552 36780 34561
rect 38292 34552 38344 34604
rect 16764 34416 16816 34468
rect 10140 34348 10192 34400
rect 11980 34348 12032 34400
rect 13912 34348 13964 34400
rect 14372 34391 14424 34400
rect 14372 34357 14381 34391
rect 14381 34357 14415 34391
rect 14415 34357 14424 34391
rect 14372 34348 14424 34357
rect 15108 34348 15160 34400
rect 17868 34348 17920 34400
rect 18512 34348 18564 34400
rect 19984 34391 20036 34400
rect 19984 34357 19993 34391
rect 19993 34357 20027 34391
rect 20027 34357 20036 34391
rect 19984 34348 20036 34357
rect 25780 34348 25832 34400
rect 28540 34484 28592 34536
rect 29000 34527 29052 34536
rect 29000 34493 29009 34527
rect 29009 34493 29043 34527
rect 29043 34493 29052 34527
rect 29000 34484 29052 34493
rect 33784 34527 33836 34536
rect 33784 34493 33793 34527
rect 33793 34493 33827 34527
rect 33827 34493 33836 34527
rect 33784 34484 33836 34493
rect 35808 34527 35860 34536
rect 35808 34493 35817 34527
rect 35817 34493 35851 34527
rect 35851 34493 35860 34527
rect 35808 34484 35860 34493
rect 28264 34416 28316 34468
rect 27344 34391 27396 34400
rect 27344 34357 27353 34391
rect 27353 34357 27387 34391
rect 27387 34357 27396 34391
rect 27344 34348 27396 34357
rect 30656 34348 30708 34400
rect 30748 34348 30800 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 3240 34144 3292 34196
rect 3792 34144 3844 34196
rect 3424 34076 3476 34128
rect 5632 34144 5684 34196
rect 6000 34144 6052 34196
rect 9864 34187 9916 34196
rect 5724 34076 5776 34128
rect 9864 34153 9873 34187
rect 9873 34153 9907 34187
rect 9907 34153 9916 34187
rect 9864 34144 9916 34153
rect 10140 34144 10192 34196
rect 11796 34144 11848 34196
rect 14464 34144 14516 34196
rect 16212 34144 16264 34196
rect 16304 34144 16356 34196
rect 17868 34144 17920 34196
rect 20996 34144 21048 34196
rect 25228 34187 25280 34196
rect 25228 34153 25237 34187
rect 25237 34153 25271 34187
rect 25271 34153 25280 34187
rect 25228 34144 25280 34153
rect 11152 34008 11204 34060
rect 5264 33872 5316 33924
rect 5816 33940 5868 33992
rect 9956 33983 10008 33992
rect 9956 33949 9965 33983
rect 9965 33949 9999 33983
rect 9999 33949 10008 33983
rect 9956 33940 10008 33949
rect 6000 33915 6052 33924
rect 6000 33881 6009 33915
rect 6009 33881 6043 33915
rect 6043 33881 6052 33915
rect 6000 33872 6052 33881
rect 7472 33915 7524 33924
rect 7472 33881 7481 33915
rect 7481 33881 7515 33915
rect 7515 33881 7524 33915
rect 7472 33872 7524 33881
rect 11796 33940 11848 33992
rect 11980 33983 12032 33992
rect 11980 33949 11989 33983
rect 11989 33949 12023 33983
rect 12023 33949 12032 33983
rect 11980 33940 12032 33949
rect 12532 33940 12584 33992
rect 13820 34008 13872 34060
rect 17040 34076 17092 34128
rect 24124 34076 24176 34128
rect 29000 34144 29052 34196
rect 29920 34187 29972 34196
rect 29920 34153 29929 34187
rect 29929 34153 29963 34187
rect 29963 34153 29972 34187
rect 29920 34144 29972 34153
rect 26976 34076 27028 34128
rect 15108 34008 15160 34060
rect 15384 34051 15436 34060
rect 15384 34017 15393 34051
rect 15393 34017 15427 34051
rect 15427 34017 15436 34051
rect 15384 34008 15436 34017
rect 16396 34008 16448 34060
rect 18604 34008 18656 34060
rect 21916 34051 21968 34060
rect 21916 34017 21925 34051
rect 21925 34017 21959 34051
rect 21959 34017 21968 34051
rect 21916 34008 21968 34017
rect 23388 34008 23440 34060
rect 27344 34008 27396 34060
rect 28724 34008 28776 34060
rect 13268 33983 13320 33992
rect 13268 33949 13277 33983
rect 13277 33949 13311 33983
rect 13311 33949 13320 33983
rect 13268 33940 13320 33949
rect 18236 33983 18288 33992
rect 11152 33872 11204 33924
rect 12624 33872 12676 33924
rect 18236 33949 18245 33983
rect 18245 33949 18279 33983
rect 18279 33949 18288 33983
rect 18236 33940 18288 33949
rect 18512 33983 18564 33992
rect 18512 33949 18521 33983
rect 18521 33949 18555 33983
rect 18555 33949 18564 33983
rect 18512 33940 18564 33949
rect 20996 33983 21048 33992
rect 20996 33949 21005 33983
rect 21005 33949 21039 33983
rect 21039 33949 21048 33983
rect 20996 33940 21048 33949
rect 24216 33940 24268 33992
rect 24676 33983 24728 33992
rect 24676 33949 24685 33983
rect 24685 33949 24719 33983
rect 24719 33949 24728 33983
rect 24676 33940 24728 33949
rect 24952 33940 25004 33992
rect 25964 33940 26016 33992
rect 26240 33983 26292 33992
rect 26240 33949 26249 33983
rect 26249 33949 26283 33983
rect 26283 33949 26292 33983
rect 26240 33940 26292 33949
rect 27712 33983 27764 33992
rect 27712 33949 27721 33983
rect 27721 33949 27755 33983
rect 27755 33949 27764 33983
rect 27712 33940 27764 33949
rect 30104 34076 30156 34128
rect 10140 33804 10192 33856
rect 11704 33804 11756 33856
rect 11888 33804 11940 33856
rect 14188 33872 14240 33924
rect 14372 33872 14424 33924
rect 15660 33915 15712 33924
rect 15660 33881 15669 33915
rect 15669 33881 15703 33915
rect 15703 33881 15712 33915
rect 15660 33872 15712 33881
rect 16948 33872 17000 33924
rect 13084 33804 13136 33856
rect 13268 33804 13320 33856
rect 15200 33804 15252 33856
rect 19340 33872 19392 33924
rect 19984 33872 20036 33924
rect 22652 33872 22704 33924
rect 26700 33872 26752 33924
rect 29920 33940 29972 33992
rect 30564 33940 30616 33992
rect 32404 34008 32456 34060
rect 37372 34051 37424 34060
rect 37372 34017 37381 34051
rect 37381 34017 37415 34051
rect 37415 34017 37424 34051
rect 37372 34008 37424 34017
rect 30932 33940 30984 33992
rect 31300 33940 31352 33992
rect 36268 33983 36320 33992
rect 36268 33949 36277 33983
rect 36277 33949 36311 33983
rect 36311 33949 36320 33983
rect 36268 33940 36320 33949
rect 27896 33872 27948 33924
rect 32312 33915 32364 33924
rect 32312 33881 32321 33915
rect 32321 33881 32355 33915
rect 32355 33881 32364 33915
rect 32312 33872 32364 33881
rect 33324 33872 33376 33924
rect 37372 33872 37424 33924
rect 18972 33804 19024 33856
rect 23480 33804 23532 33856
rect 24400 33847 24452 33856
rect 24400 33813 24409 33847
rect 24409 33813 24443 33847
rect 24443 33813 24452 33847
rect 24400 33804 24452 33813
rect 26332 33804 26384 33856
rect 27528 33847 27580 33856
rect 27528 33813 27537 33847
rect 27537 33813 27571 33847
rect 27571 33813 27580 33847
rect 27528 33804 27580 33813
rect 30012 33804 30064 33856
rect 32128 33804 32180 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 5356 33600 5408 33652
rect 11060 33532 11112 33584
rect 2964 33464 3016 33516
rect 3608 33507 3660 33516
rect 3608 33473 3617 33507
rect 3617 33473 3651 33507
rect 3651 33473 3660 33507
rect 3608 33464 3660 33473
rect 5816 33464 5868 33516
rect 6736 33464 6788 33516
rect 10232 33464 10284 33516
rect 5356 33439 5408 33448
rect 5356 33405 5365 33439
rect 5365 33405 5399 33439
rect 5399 33405 5408 33439
rect 5356 33396 5408 33405
rect 10876 33464 10928 33516
rect 3424 33328 3476 33380
rect 10140 33328 10192 33380
rect 11152 33396 11204 33448
rect 10692 33328 10744 33380
rect 8392 33260 8444 33312
rect 9128 33303 9180 33312
rect 9128 33269 9137 33303
rect 9137 33269 9171 33303
rect 9171 33269 9180 33303
rect 9128 33260 9180 33269
rect 10324 33303 10376 33312
rect 10324 33269 10333 33303
rect 10333 33269 10367 33303
rect 10367 33269 10376 33303
rect 10324 33260 10376 33269
rect 10784 33303 10836 33312
rect 10784 33269 10793 33303
rect 10793 33269 10827 33303
rect 10827 33269 10836 33303
rect 10784 33260 10836 33269
rect 14556 33600 14608 33652
rect 16488 33600 16540 33652
rect 17040 33600 17092 33652
rect 18236 33600 18288 33652
rect 22468 33600 22520 33652
rect 24400 33600 24452 33652
rect 24952 33643 25004 33652
rect 24952 33609 24961 33643
rect 24961 33609 24995 33643
rect 24995 33609 25004 33643
rect 24952 33600 25004 33609
rect 25872 33600 25924 33652
rect 26240 33600 26292 33652
rect 33324 33600 33376 33652
rect 37372 33643 37424 33652
rect 37372 33609 37381 33643
rect 37381 33609 37415 33643
rect 37415 33609 37424 33643
rect 37372 33600 37424 33609
rect 11796 33532 11848 33584
rect 12808 33532 12860 33584
rect 15200 33532 15252 33584
rect 15292 33532 15344 33584
rect 17408 33532 17460 33584
rect 18420 33532 18472 33584
rect 20720 33532 20772 33584
rect 20996 33532 21048 33584
rect 23388 33575 23440 33584
rect 23388 33541 23397 33575
rect 23397 33541 23431 33575
rect 23431 33541 23440 33575
rect 23388 33532 23440 33541
rect 12348 33396 12400 33448
rect 12900 33439 12952 33448
rect 12900 33405 12909 33439
rect 12909 33405 12943 33439
rect 12943 33405 12952 33439
rect 12900 33396 12952 33405
rect 13360 33396 13412 33448
rect 11520 33371 11572 33380
rect 11520 33337 11529 33371
rect 11529 33337 11563 33371
rect 11563 33337 11572 33371
rect 11520 33328 11572 33337
rect 14280 33396 14332 33448
rect 15292 33439 15344 33448
rect 15292 33405 15301 33439
rect 15301 33405 15335 33439
rect 15335 33405 15344 33439
rect 15292 33396 15344 33405
rect 24032 33464 24084 33516
rect 17592 33439 17644 33448
rect 17592 33405 17601 33439
rect 17601 33405 17635 33439
rect 17635 33405 17644 33439
rect 17592 33396 17644 33405
rect 18696 33439 18748 33448
rect 18696 33405 18705 33439
rect 18705 33405 18739 33439
rect 18739 33405 18748 33439
rect 18696 33396 18748 33405
rect 18972 33439 19024 33448
rect 18972 33405 18981 33439
rect 18981 33405 19015 33439
rect 19015 33405 19024 33439
rect 19524 33439 19576 33448
rect 18972 33396 19024 33405
rect 19524 33405 19533 33439
rect 19533 33405 19567 33439
rect 19567 33405 19576 33439
rect 19524 33396 19576 33405
rect 20904 33396 20956 33448
rect 23480 33439 23532 33448
rect 23480 33405 23489 33439
rect 23489 33405 23523 33439
rect 23523 33405 23532 33439
rect 23480 33396 23532 33405
rect 25228 33532 25280 33584
rect 30012 33532 30064 33584
rect 30196 33532 30248 33584
rect 25044 33464 25096 33516
rect 25596 33507 25648 33516
rect 25596 33473 25605 33507
rect 25605 33473 25639 33507
rect 25639 33473 25648 33507
rect 25596 33464 25648 33473
rect 26976 33507 27028 33516
rect 26976 33473 26985 33507
rect 26985 33473 27019 33507
rect 27019 33473 27028 33507
rect 26976 33464 27028 33473
rect 27896 33507 27948 33516
rect 27896 33473 27905 33507
rect 27905 33473 27939 33507
rect 27939 33473 27948 33507
rect 27896 33464 27948 33473
rect 28172 33464 28224 33516
rect 32128 33507 32180 33516
rect 32128 33473 32137 33507
rect 32137 33473 32171 33507
rect 32171 33473 32180 33507
rect 32128 33464 32180 33473
rect 32404 33464 32456 33516
rect 34704 33464 34756 33516
rect 36268 33464 36320 33516
rect 38108 33507 38160 33516
rect 24584 33439 24636 33448
rect 24584 33405 24593 33439
rect 24593 33405 24627 33439
rect 24627 33405 24636 33439
rect 24584 33396 24636 33405
rect 16764 33260 16816 33312
rect 18604 33260 18656 33312
rect 23572 33260 23624 33312
rect 24400 33260 24452 33312
rect 24860 33396 24912 33448
rect 25412 33439 25464 33448
rect 25412 33405 25421 33439
rect 25421 33405 25455 33439
rect 25455 33405 25464 33439
rect 25412 33396 25464 33405
rect 27804 33439 27856 33448
rect 27804 33405 27813 33439
rect 27813 33405 27847 33439
rect 27847 33405 27856 33439
rect 27804 33396 27856 33405
rect 27988 33439 28040 33448
rect 27988 33405 27997 33439
rect 27997 33405 28031 33439
rect 28031 33405 28040 33439
rect 27988 33396 28040 33405
rect 30932 33396 30984 33448
rect 31024 33396 31076 33448
rect 38108 33473 38117 33507
rect 38117 33473 38151 33507
rect 38151 33473 38160 33507
rect 38108 33464 38160 33473
rect 37556 33396 37608 33448
rect 24952 33260 25004 33312
rect 27068 33303 27120 33312
rect 27068 33269 27077 33303
rect 27077 33269 27111 33303
rect 27111 33269 27120 33303
rect 27068 33260 27120 33269
rect 29000 33303 29052 33312
rect 29000 33269 29009 33303
rect 29009 33269 29043 33303
rect 29043 33269 29052 33303
rect 29000 33260 29052 33269
rect 30840 33260 30892 33312
rect 31760 33260 31812 33312
rect 32036 33260 32088 33312
rect 32956 33260 33008 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 10324 33056 10376 33108
rect 11244 33056 11296 33108
rect 10876 32988 10928 33040
rect 5816 32895 5868 32904
rect 5816 32861 5825 32895
rect 5825 32861 5859 32895
rect 5859 32861 5868 32895
rect 5816 32852 5868 32861
rect 4712 32784 4764 32836
rect 8484 32920 8536 32972
rect 11520 32920 11572 32972
rect 7748 32895 7800 32904
rect 7748 32861 7757 32895
rect 7757 32861 7791 32895
rect 7791 32861 7800 32895
rect 7748 32852 7800 32861
rect 7840 32895 7892 32904
rect 7840 32861 7849 32895
rect 7849 32861 7883 32895
rect 7883 32861 7892 32895
rect 7840 32852 7892 32861
rect 11612 32895 11664 32904
rect 7380 32716 7432 32768
rect 9128 32784 9180 32836
rect 10416 32827 10468 32836
rect 10416 32793 10425 32827
rect 10425 32793 10459 32827
rect 10459 32793 10468 32827
rect 10416 32784 10468 32793
rect 9772 32716 9824 32768
rect 10048 32716 10100 32768
rect 11612 32861 11621 32895
rect 11621 32861 11655 32895
rect 11655 32861 11664 32895
rect 11612 32852 11664 32861
rect 11888 32852 11940 32904
rect 12900 33056 12952 33108
rect 14648 33056 14700 33108
rect 18420 33099 18472 33108
rect 14280 32988 14332 33040
rect 18420 33065 18429 33099
rect 18429 33065 18463 33099
rect 18463 33065 18472 33099
rect 18420 33056 18472 33065
rect 20720 33099 20772 33108
rect 20720 33065 20729 33099
rect 20729 33065 20763 33099
rect 20763 33065 20772 33099
rect 20720 33056 20772 33065
rect 22652 33056 22704 33108
rect 24584 33056 24636 33108
rect 15384 32920 15436 32972
rect 18236 32920 18288 32972
rect 13084 32895 13136 32904
rect 13084 32861 13093 32895
rect 13093 32861 13127 32895
rect 13127 32861 13136 32895
rect 13084 32852 13136 32861
rect 14004 32852 14056 32904
rect 15292 32852 15344 32904
rect 18420 32852 18472 32904
rect 18972 32852 19024 32904
rect 19156 32852 19208 32904
rect 19524 32895 19576 32904
rect 19524 32861 19533 32895
rect 19533 32861 19567 32895
rect 19567 32861 19576 32895
rect 19524 32852 19576 32861
rect 20904 32988 20956 33040
rect 24400 32988 24452 33040
rect 28172 33056 28224 33108
rect 28540 33056 28592 33108
rect 30196 33099 30248 33108
rect 30196 33065 30205 33099
rect 30205 33065 30239 33099
rect 30239 33065 30248 33099
rect 30196 33056 30248 33065
rect 30656 33099 30708 33108
rect 30656 33065 30665 33099
rect 30665 33065 30699 33099
rect 30699 33065 30708 33099
rect 30656 33056 30708 33065
rect 30748 33056 30800 33108
rect 31024 32988 31076 33040
rect 26056 32963 26108 32972
rect 20076 32852 20128 32904
rect 20812 32895 20864 32904
rect 20812 32861 20821 32895
rect 20821 32861 20855 32895
rect 20855 32861 20864 32895
rect 20812 32852 20864 32861
rect 21456 32852 21508 32904
rect 14648 32784 14700 32836
rect 15200 32784 15252 32836
rect 17040 32784 17092 32836
rect 18604 32784 18656 32836
rect 21732 32827 21784 32836
rect 21732 32793 21741 32827
rect 21741 32793 21775 32827
rect 21775 32793 21784 32827
rect 26056 32929 26065 32963
rect 26065 32929 26099 32963
rect 26099 32929 26108 32963
rect 26056 32920 26108 32929
rect 26332 32963 26384 32972
rect 26332 32929 26341 32963
rect 26341 32929 26375 32963
rect 26375 32929 26384 32963
rect 26332 32920 26384 32929
rect 26424 32920 26476 32972
rect 23388 32852 23440 32904
rect 23480 32852 23532 32904
rect 24492 32852 24544 32904
rect 27896 32920 27948 32972
rect 30472 32920 30524 32972
rect 28540 32852 28592 32904
rect 21732 32784 21784 32793
rect 24308 32784 24360 32836
rect 25044 32784 25096 32836
rect 11796 32716 11848 32768
rect 14188 32759 14240 32768
rect 14188 32725 14197 32759
rect 14197 32725 14231 32759
rect 14231 32725 14240 32759
rect 14188 32716 14240 32725
rect 16488 32716 16540 32768
rect 18328 32716 18380 32768
rect 22928 32716 22980 32768
rect 23572 32759 23624 32768
rect 23572 32725 23599 32759
rect 23599 32725 23624 32759
rect 23572 32716 23624 32725
rect 24216 32716 24268 32768
rect 24952 32716 25004 32768
rect 25504 32759 25556 32768
rect 25504 32725 25513 32759
rect 25513 32725 25547 32759
rect 25547 32725 25556 32759
rect 25504 32716 25556 32725
rect 26424 32716 26476 32768
rect 27068 32784 27120 32836
rect 28724 32895 28776 32904
rect 28724 32861 28733 32895
rect 28733 32861 28767 32895
rect 28767 32861 28776 32895
rect 28724 32852 28776 32861
rect 29000 32852 29052 32904
rect 29828 32852 29880 32904
rect 30104 32852 30156 32904
rect 30840 32895 30892 32904
rect 30840 32861 30849 32895
rect 30849 32861 30883 32895
rect 30883 32861 30892 32895
rect 30840 32852 30892 32861
rect 31576 33056 31628 33108
rect 31760 33099 31812 33108
rect 31760 33065 31769 33099
rect 31769 33065 31803 33099
rect 31803 33065 31812 33099
rect 31760 33056 31812 33065
rect 31852 33056 31904 33108
rect 33600 33056 33652 33108
rect 31944 32963 31996 32972
rect 31944 32929 31953 32963
rect 31953 32929 31987 32963
rect 31987 32929 31996 32963
rect 31944 32920 31996 32929
rect 32496 32920 32548 32972
rect 31024 32861 31033 32882
rect 31033 32861 31067 32882
rect 31067 32861 31076 32882
rect 31024 32830 31076 32861
rect 31300 32895 31352 32904
rect 31300 32861 31309 32895
rect 31309 32861 31343 32895
rect 31343 32861 31352 32895
rect 32036 32895 32088 32904
rect 31300 32852 31352 32861
rect 32036 32861 32045 32895
rect 32045 32861 32079 32895
rect 32079 32861 32088 32895
rect 32036 32852 32088 32861
rect 32772 32895 32824 32904
rect 28448 32716 28500 32768
rect 31576 32784 31628 32836
rect 32772 32861 32781 32895
rect 32781 32861 32815 32895
rect 32815 32861 32824 32895
rect 32772 32852 32824 32861
rect 34704 32895 34756 32904
rect 34704 32861 34713 32895
rect 34713 32861 34747 32895
rect 34747 32861 34756 32895
rect 34704 32852 34756 32861
rect 36268 32895 36320 32904
rect 36268 32861 36277 32895
rect 36277 32861 36311 32895
rect 36311 32861 36320 32895
rect 36268 32852 36320 32861
rect 32956 32827 33008 32836
rect 32956 32793 32965 32827
rect 32965 32793 32999 32827
rect 32999 32793 33008 32827
rect 32956 32784 33008 32793
rect 33692 32784 33744 32836
rect 37648 32784 37700 32836
rect 38108 32827 38160 32836
rect 38108 32793 38117 32827
rect 38117 32793 38151 32827
rect 38151 32793 38160 32827
rect 38108 32784 38160 32793
rect 31760 32716 31812 32768
rect 32404 32716 32456 32768
rect 34060 32716 34112 32768
rect 34796 32759 34848 32768
rect 34796 32725 34805 32759
rect 34805 32725 34839 32759
rect 34839 32725 34848 32759
rect 34796 32716 34848 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 6736 32444 6788 32496
rect 6828 32419 6880 32428
rect 6828 32385 6837 32419
rect 6837 32385 6871 32419
rect 6871 32385 6880 32419
rect 6828 32376 6880 32385
rect 7012 32419 7064 32428
rect 7012 32385 7021 32419
rect 7021 32385 7055 32419
rect 7055 32385 7064 32419
rect 7012 32376 7064 32385
rect 6552 32308 6604 32360
rect 8484 32512 8536 32564
rect 8392 32444 8444 32496
rect 10416 32512 10468 32564
rect 12808 32512 12860 32564
rect 13084 32555 13136 32564
rect 13084 32521 13093 32555
rect 13093 32521 13127 32555
rect 13127 32521 13136 32555
rect 13084 32512 13136 32521
rect 15200 32555 15252 32564
rect 15200 32521 15209 32555
rect 15209 32521 15243 32555
rect 15243 32521 15252 32555
rect 15200 32512 15252 32521
rect 15384 32512 15436 32564
rect 19248 32512 19300 32564
rect 20996 32512 21048 32564
rect 11060 32444 11112 32496
rect 12992 32444 13044 32496
rect 15292 32444 15344 32496
rect 15476 32487 15528 32496
rect 15476 32453 15485 32487
rect 15485 32453 15519 32487
rect 15519 32453 15528 32487
rect 15476 32444 15528 32453
rect 16488 32444 16540 32496
rect 10048 32376 10100 32428
rect 10416 32376 10468 32428
rect 11704 32419 11756 32428
rect 11704 32385 11713 32419
rect 11713 32385 11747 32419
rect 11747 32385 11756 32419
rect 11704 32376 11756 32385
rect 11796 32419 11848 32428
rect 11796 32385 11805 32419
rect 11805 32385 11839 32419
rect 11839 32385 11848 32419
rect 11796 32376 11848 32385
rect 12256 32376 12308 32428
rect 15384 32419 15436 32428
rect 15384 32385 15393 32419
rect 15393 32385 15427 32419
rect 15427 32385 15436 32419
rect 15384 32376 15436 32385
rect 15568 32419 15620 32428
rect 15568 32385 15577 32419
rect 15577 32385 15611 32419
rect 15611 32385 15620 32419
rect 15568 32376 15620 32385
rect 19432 32444 19484 32496
rect 25964 32512 26016 32564
rect 26976 32512 27028 32564
rect 27804 32555 27856 32564
rect 27804 32521 27831 32555
rect 27831 32521 27856 32555
rect 27804 32512 27856 32521
rect 28908 32512 28960 32564
rect 30104 32555 30156 32564
rect 30104 32521 30113 32555
rect 30113 32521 30147 32555
rect 30147 32521 30156 32555
rect 30104 32512 30156 32521
rect 30656 32512 30708 32564
rect 32036 32512 32088 32564
rect 32312 32512 32364 32564
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 3240 32172 3292 32224
rect 5724 32215 5776 32224
rect 5724 32181 5733 32215
rect 5733 32181 5767 32215
rect 5767 32181 5776 32215
rect 5724 32172 5776 32181
rect 8392 32172 8444 32224
rect 10876 32308 10928 32360
rect 12164 32351 12216 32360
rect 10416 32172 10468 32224
rect 12164 32317 12173 32351
rect 12173 32317 12207 32351
rect 12207 32317 12216 32351
rect 12164 32308 12216 32317
rect 11060 32240 11112 32292
rect 17224 32376 17276 32428
rect 18696 32376 18748 32428
rect 16856 32308 16908 32360
rect 19156 32376 19208 32428
rect 21088 32419 21140 32428
rect 19064 32308 19116 32360
rect 19340 32308 19392 32360
rect 11612 32172 11664 32224
rect 13360 32172 13412 32224
rect 16764 32240 16816 32292
rect 21088 32385 21097 32419
rect 21097 32385 21131 32419
rect 21131 32385 21140 32419
rect 21088 32376 21140 32385
rect 22560 32444 22612 32496
rect 24032 32444 24084 32496
rect 25504 32444 25556 32496
rect 24584 32376 24636 32428
rect 25872 32444 25924 32496
rect 26424 32444 26476 32496
rect 26056 32419 26108 32428
rect 26056 32385 26065 32419
rect 26065 32385 26099 32419
rect 26099 32385 26108 32419
rect 26056 32376 26108 32385
rect 27068 32376 27120 32428
rect 28172 32444 28224 32496
rect 29184 32444 29236 32496
rect 29736 32487 29788 32496
rect 29736 32453 29745 32487
rect 29745 32453 29779 32487
rect 29779 32453 29788 32487
rect 29736 32444 29788 32453
rect 29828 32444 29880 32496
rect 31116 32487 31168 32496
rect 31116 32453 31125 32487
rect 31125 32453 31159 32487
rect 31159 32453 31168 32487
rect 31116 32444 31168 32453
rect 23572 32351 23624 32360
rect 23572 32317 23581 32351
rect 23581 32317 23615 32351
rect 23615 32317 23624 32351
rect 23572 32308 23624 32317
rect 24216 32351 24268 32360
rect 24216 32317 24225 32351
rect 24225 32317 24259 32351
rect 24259 32317 24268 32351
rect 24216 32308 24268 32317
rect 24308 32351 24360 32360
rect 24308 32317 24317 32351
rect 24317 32317 24351 32351
rect 24351 32317 24360 32351
rect 24492 32351 24544 32360
rect 24308 32308 24360 32317
rect 24492 32317 24501 32351
rect 24501 32317 24535 32351
rect 24535 32317 24544 32351
rect 24492 32308 24544 32317
rect 25228 32308 25280 32360
rect 25688 32308 25740 32360
rect 30196 32376 30248 32428
rect 30288 32376 30340 32428
rect 31668 32444 31720 32496
rect 31852 32444 31904 32496
rect 34704 32512 34756 32564
rect 37648 32555 37700 32564
rect 37648 32521 37657 32555
rect 37657 32521 37691 32555
rect 37691 32521 37700 32555
rect 37648 32512 37700 32521
rect 25596 32240 25648 32292
rect 27712 32240 27764 32292
rect 28448 32283 28500 32292
rect 28448 32249 28457 32283
rect 28457 32249 28491 32283
rect 28491 32249 28500 32283
rect 31760 32308 31812 32360
rect 32864 32444 32916 32496
rect 32404 32419 32456 32428
rect 32404 32385 32413 32419
rect 32413 32385 32447 32419
rect 32447 32385 32456 32419
rect 32404 32376 32456 32385
rect 32312 32308 32364 32360
rect 32956 32376 33008 32428
rect 34796 32376 34848 32428
rect 36268 32376 36320 32428
rect 37924 32376 37976 32428
rect 33232 32308 33284 32360
rect 33416 32351 33468 32360
rect 33416 32317 33425 32351
rect 33425 32317 33459 32351
rect 33459 32317 33468 32351
rect 33416 32308 33468 32317
rect 34152 32308 34204 32360
rect 28448 32240 28500 32249
rect 18696 32172 18748 32224
rect 18880 32172 18932 32224
rect 19340 32172 19392 32224
rect 22100 32172 22152 32224
rect 27344 32172 27396 32224
rect 27988 32172 28040 32224
rect 28632 32215 28684 32224
rect 28632 32181 28641 32215
rect 28641 32181 28675 32215
rect 28675 32181 28684 32215
rect 28632 32172 28684 32181
rect 28816 32172 28868 32224
rect 30748 32240 30800 32292
rect 31944 32240 31996 32292
rect 36268 32172 36320 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 7656 31968 7708 32020
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 3240 31875 3292 31884
rect 3240 31841 3249 31875
rect 3249 31841 3283 31875
rect 3283 31841 3292 31875
rect 3240 31832 3292 31841
rect 7840 31900 7892 31952
rect 11704 31968 11756 32020
rect 11796 31968 11848 32020
rect 13176 31968 13228 32020
rect 16764 31968 16816 32020
rect 18052 31968 18104 32020
rect 7288 31875 7340 31884
rect 7288 31841 7297 31875
rect 7297 31841 7331 31875
rect 7331 31841 7340 31875
rect 11060 31900 11112 31952
rect 15292 31900 15344 31952
rect 17224 31943 17276 31952
rect 17224 31909 17233 31943
rect 17233 31909 17267 31943
rect 17267 31909 17276 31943
rect 17224 31900 17276 31909
rect 7288 31832 7340 31841
rect 11704 31832 11756 31884
rect 6552 31807 6604 31816
rect 6552 31773 6561 31807
rect 6561 31773 6595 31807
rect 6595 31773 6604 31807
rect 6552 31764 6604 31773
rect 7380 31807 7432 31816
rect 7380 31773 7389 31807
rect 7389 31773 7423 31807
rect 7423 31773 7432 31807
rect 7656 31807 7708 31816
rect 7380 31764 7432 31773
rect 7656 31773 7665 31807
rect 7665 31773 7699 31807
rect 7699 31773 7708 31807
rect 7656 31764 7708 31773
rect 7840 31764 7892 31816
rect 3056 31739 3108 31748
rect 3056 31705 3065 31739
rect 3065 31705 3099 31739
rect 3099 31705 3108 31739
rect 3056 31696 3108 31705
rect 5724 31696 5776 31748
rect 7380 31628 7432 31680
rect 8300 31764 8352 31816
rect 9864 31764 9916 31816
rect 10232 31807 10284 31816
rect 10232 31773 10241 31807
rect 10241 31773 10275 31807
rect 10275 31773 10284 31807
rect 10232 31764 10284 31773
rect 11060 31807 11112 31816
rect 11060 31773 11069 31807
rect 11069 31773 11103 31807
rect 11103 31773 11112 31807
rect 11060 31764 11112 31773
rect 10416 31739 10468 31748
rect 10416 31705 10425 31739
rect 10425 31705 10459 31739
rect 10459 31705 10468 31739
rect 10416 31696 10468 31705
rect 12164 31764 12216 31816
rect 14004 31832 14056 31884
rect 13544 31764 13596 31816
rect 15016 31764 15068 31816
rect 15200 31764 15252 31816
rect 16856 31832 16908 31884
rect 18972 31832 19024 31884
rect 15660 31764 15712 31816
rect 16304 31807 16356 31816
rect 16304 31773 16313 31807
rect 16313 31773 16347 31807
rect 16347 31773 16356 31807
rect 16304 31764 16356 31773
rect 16488 31807 16540 31816
rect 16488 31773 16497 31807
rect 16497 31773 16531 31807
rect 16531 31773 16540 31807
rect 16488 31764 16540 31773
rect 17684 31807 17736 31816
rect 17684 31773 17693 31807
rect 17693 31773 17727 31807
rect 17727 31773 17736 31807
rect 17684 31764 17736 31773
rect 17868 31807 17920 31816
rect 17868 31773 17877 31807
rect 17877 31773 17911 31807
rect 17911 31773 17920 31807
rect 17868 31764 17920 31773
rect 13268 31696 13320 31748
rect 18512 31739 18564 31748
rect 18512 31705 18539 31739
rect 18539 31705 18564 31739
rect 18512 31696 18564 31705
rect 18788 31696 18840 31748
rect 21088 31968 21140 32020
rect 24124 31968 24176 32020
rect 24400 31968 24452 32020
rect 29092 31968 29144 32020
rect 30288 31968 30340 32020
rect 19248 31875 19300 31884
rect 19248 31841 19257 31875
rect 19257 31841 19291 31875
rect 19291 31841 19300 31875
rect 19248 31832 19300 31841
rect 28172 31900 28224 31952
rect 22836 31832 22888 31884
rect 23572 31832 23624 31884
rect 20628 31764 20680 31816
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22100 31807 22152 31816
rect 22100 31773 22109 31807
rect 22109 31773 22143 31807
rect 22143 31773 22152 31807
rect 22100 31764 22152 31773
rect 23388 31764 23440 31816
rect 24308 31764 24360 31816
rect 25412 31807 25464 31816
rect 25412 31773 25421 31807
rect 25421 31773 25455 31807
rect 25455 31773 25464 31807
rect 25412 31764 25464 31773
rect 26056 31764 26108 31816
rect 19432 31696 19484 31748
rect 22928 31739 22980 31748
rect 22928 31705 22937 31739
rect 22937 31705 22971 31739
rect 22971 31705 22980 31739
rect 22928 31696 22980 31705
rect 24400 31739 24452 31748
rect 24400 31705 24409 31739
rect 24409 31705 24443 31739
rect 24443 31705 24452 31739
rect 24400 31696 24452 31705
rect 24584 31739 24636 31748
rect 24584 31705 24593 31739
rect 24593 31705 24627 31739
rect 24627 31705 24636 31739
rect 24584 31696 24636 31705
rect 25044 31696 25096 31748
rect 18144 31628 18196 31680
rect 25872 31628 25924 31680
rect 27528 31832 27580 31884
rect 27988 31832 28040 31884
rect 29184 31900 29236 31952
rect 31576 31968 31628 32020
rect 34612 31968 34664 32020
rect 27620 31764 27672 31816
rect 29828 31832 29880 31884
rect 30288 31832 30340 31884
rect 30840 31832 30892 31884
rect 32128 31900 32180 31952
rect 33692 31900 33744 31952
rect 29920 31764 29972 31816
rect 26792 31628 26844 31680
rect 27804 31696 27856 31748
rect 30472 31696 30524 31748
rect 31116 31764 31168 31816
rect 32956 31832 33008 31884
rect 33232 31832 33284 31884
rect 31668 31807 31720 31816
rect 31668 31773 31677 31807
rect 31677 31773 31711 31807
rect 31711 31773 31720 31807
rect 31668 31764 31720 31773
rect 31944 31764 31996 31816
rect 32496 31764 32548 31816
rect 34060 31832 34112 31884
rect 34152 31875 34204 31884
rect 34152 31841 34161 31875
rect 34161 31841 34195 31875
rect 34195 31841 34204 31875
rect 34704 31875 34756 31884
rect 34152 31832 34204 31841
rect 34704 31841 34713 31875
rect 34713 31841 34747 31875
rect 34747 31841 34756 31875
rect 34704 31832 34756 31841
rect 36268 31875 36320 31884
rect 36268 31841 36277 31875
rect 36277 31841 36311 31875
rect 36311 31841 36320 31875
rect 36268 31832 36320 31841
rect 38108 31807 38160 31816
rect 38108 31773 38117 31807
rect 38117 31773 38151 31807
rect 38151 31773 38160 31807
rect 38108 31764 38160 31773
rect 31576 31696 31628 31748
rect 33784 31739 33836 31748
rect 33784 31705 33793 31739
rect 33793 31705 33827 31739
rect 33827 31705 33836 31739
rect 33784 31696 33836 31705
rect 33876 31739 33928 31748
rect 33876 31705 33885 31739
rect 33885 31705 33919 31739
rect 33919 31705 33928 31739
rect 36452 31739 36504 31748
rect 33876 31696 33928 31705
rect 36452 31705 36461 31739
rect 36461 31705 36495 31739
rect 36495 31705 36504 31739
rect 36452 31696 36504 31705
rect 28356 31628 28408 31680
rect 29920 31628 29972 31680
rect 30012 31628 30064 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 3056 31424 3108 31476
rect 6828 31424 6880 31476
rect 7748 31424 7800 31476
rect 2320 31288 2372 31340
rect 7288 31356 7340 31408
rect 5908 31288 5960 31340
rect 7748 31331 7800 31340
rect 7748 31297 7757 31331
rect 7757 31297 7791 31331
rect 7791 31297 7800 31331
rect 7748 31288 7800 31297
rect 9864 31424 9916 31476
rect 11060 31424 11112 31476
rect 16028 31424 16080 31476
rect 16396 31424 16448 31476
rect 17684 31467 17736 31476
rect 17684 31433 17693 31467
rect 17693 31433 17727 31467
rect 17727 31433 17736 31467
rect 17684 31424 17736 31433
rect 18144 31424 18196 31476
rect 19064 31424 19116 31476
rect 19432 31424 19484 31476
rect 20628 31467 20680 31476
rect 20628 31433 20637 31467
rect 20637 31433 20671 31467
rect 20671 31433 20680 31467
rect 20628 31424 20680 31433
rect 22560 31424 22612 31476
rect 22836 31424 22888 31476
rect 24216 31467 24268 31476
rect 24216 31433 24225 31467
rect 24225 31433 24259 31467
rect 24259 31433 24268 31467
rect 24216 31424 24268 31433
rect 24308 31424 24360 31476
rect 25320 31424 25372 31476
rect 27804 31424 27856 31476
rect 7932 31288 7984 31340
rect 8208 31288 8260 31340
rect 9496 31356 9548 31408
rect 7288 31220 7340 31272
rect 7472 31195 7524 31204
rect 7472 31161 7481 31195
rect 7481 31161 7515 31195
rect 7515 31161 7524 31195
rect 7472 31152 7524 31161
rect 5080 31127 5132 31136
rect 5080 31093 5089 31127
rect 5089 31093 5123 31127
rect 5123 31093 5132 31127
rect 5080 31084 5132 31093
rect 5172 31084 5224 31136
rect 6736 31084 6788 31136
rect 10048 31288 10100 31340
rect 10232 31288 10284 31340
rect 10876 31356 10928 31408
rect 11520 31399 11572 31408
rect 11520 31365 11529 31399
rect 11529 31365 11563 31399
rect 11563 31365 11572 31399
rect 11520 31356 11572 31365
rect 14280 31356 14332 31408
rect 16488 31356 16540 31408
rect 18420 31356 18472 31408
rect 12348 31331 12400 31340
rect 12348 31297 12357 31331
rect 12357 31297 12391 31331
rect 12391 31297 12400 31331
rect 12348 31288 12400 31297
rect 15016 31288 15068 31340
rect 15660 31331 15712 31340
rect 15660 31297 15669 31331
rect 15669 31297 15703 31331
rect 15703 31297 15712 31331
rect 15660 31288 15712 31297
rect 16396 31288 16448 31340
rect 16580 31288 16632 31340
rect 17408 31288 17460 31340
rect 18052 31331 18104 31340
rect 11612 31220 11664 31272
rect 12716 31220 12768 31272
rect 12992 31220 13044 31272
rect 18052 31297 18061 31331
rect 18061 31297 18095 31331
rect 18095 31297 18104 31331
rect 18052 31288 18104 31297
rect 18144 31331 18196 31340
rect 18144 31297 18153 31331
rect 18153 31297 18187 31331
rect 18187 31297 18196 31331
rect 18144 31288 18196 31297
rect 18512 31288 18564 31340
rect 18420 31220 18472 31272
rect 18788 31288 18840 31340
rect 18972 31331 19024 31340
rect 18972 31297 18981 31331
rect 18981 31297 19015 31331
rect 19015 31297 19024 31331
rect 18972 31288 19024 31297
rect 19064 31331 19116 31340
rect 19064 31297 19073 31331
rect 19073 31297 19107 31331
rect 19107 31297 19116 31331
rect 19064 31288 19116 31297
rect 19984 31288 20036 31340
rect 20168 31288 20220 31340
rect 20720 31331 20772 31340
rect 20720 31297 20729 31331
rect 20729 31297 20763 31331
rect 20763 31297 20772 31331
rect 20720 31288 20772 31297
rect 23388 31356 23440 31408
rect 24584 31399 24636 31408
rect 24584 31365 24593 31399
rect 24593 31365 24627 31399
rect 24627 31365 24636 31399
rect 24584 31356 24636 31365
rect 25412 31356 25464 31408
rect 27068 31356 27120 31408
rect 25044 31331 25096 31340
rect 25044 31297 25053 31331
rect 25053 31297 25087 31331
rect 25087 31297 25096 31331
rect 25044 31288 25096 31297
rect 26056 31288 26108 31340
rect 26516 31288 26568 31340
rect 26608 31288 26660 31340
rect 28356 31331 28408 31340
rect 28356 31297 28365 31331
rect 28365 31297 28399 31331
rect 28399 31297 28408 31331
rect 28356 31288 28408 31297
rect 18696 31263 18748 31272
rect 18696 31229 18705 31263
rect 18705 31229 18739 31263
rect 18739 31229 18748 31263
rect 18696 31220 18748 31229
rect 20904 31220 20956 31272
rect 23664 31220 23716 31272
rect 24400 31220 24452 31272
rect 28724 31220 28776 31272
rect 8300 31084 8352 31136
rect 9588 31127 9640 31136
rect 9588 31093 9597 31127
rect 9597 31093 9631 31127
rect 9631 31093 9640 31127
rect 9588 31084 9640 31093
rect 14372 31152 14424 31204
rect 14556 31195 14608 31204
rect 14556 31161 14565 31195
rect 14565 31161 14599 31195
rect 14599 31161 14608 31195
rect 14556 31152 14608 31161
rect 16120 31152 16172 31204
rect 22008 31152 22060 31204
rect 25872 31152 25924 31204
rect 26148 31195 26200 31204
rect 26148 31161 26157 31195
rect 26157 31161 26191 31195
rect 26191 31161 26200 31195
rect 26148 31152 26200 31161
rect 29920 31356 29972 31408
rect 30380 31424 30432 31476
rect 30656 31356 30708 31408
rect 30656 31263 30708 31272
rect 30656 31229 30665 31263
rect 30665 31229 30699 31263
rect 30699 31229 30708 31263
rect 30656 31220 30708 31229
rect 30932 31263 30984 31272
rect 30932 31229 30941 31263
rect 30941 31229 30975 31263
rect 30975 31229 30984 31263
rect 30932 31220 30984 31229
rect 31760 31424 31812 31476
rect 32864 31424 32916 31476
rect 33876 31467 33928 31476
rect 33876 31433 33885 31467
rect 33885 31433 33919 31467
rect 33919 31433 33928 31467
rect 33876 31424 33928 31433
rect 36452 31424 36504 31476
rect 32496 31356 32548 31408
rect 31484 31288 31536 31340
rect 33692 31288 33744 31340
rect 34612 31331 34664 31340
rect 34612 31297 34621 31331
rect 34621 31297 34655 31331
rect 34655 31297 34664 31331
rect 34612 31288 34664 31297
rect 36912 31288 36964 31340
rect 37924 31288 37976 31340
rect 10140 31084 10192 31136
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 11704 31127 11756 31136
rect 11704 31093 11713 31127
rect 11713 31093 11747 31127
rect 11747 31093 11756 31127
rect 11704 31084 11756 31093
rect 12164 31084 12216 31136
rect 12348 31084 12400 31136
rect 13360 31084 13412 31136
rect 15476 31084 15528 31136
rect 22560 31084 22612 31136
rect 27160 31084 27212 31136
rect 31116 31152 31168 31204
rect 32312 31152 32364 31204
rect 28540 31127 28592 31136
rect 28540 31093 28549 31127
rect 28549 31093 28583 31127
rect 28583 31093 28592 31127
rect 28540 31084 28592 31093
rect 29184 31127 29236 31136
rect 29184 31093 29193 31127
rect 29193 31093 29227 31127
rect 29227 31093 29236 31127
rect 29184 31084 29236 31093
rect 29920 31084 29972 31136
rect 33048 31084 33100 31136
rect 35440 31127 35492 31136
rect 35440 31093 35449 31127
rect 35449 31093 35483 31127
rect 35483 31093 35492 31127
rect 35440 31084 35492 31093
rect 36084 31127 36136 31136
rect 36084 31093 36093 31127
rect 36093 31093 36127 31127
rect 36127 31093 36136 31127
rect 36084 31084 36136 31093
rect 36452 31084 36504 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7748 30880 7800 30932
rect 9496 30923 9548 30932
rect 9496 30889 9505 30923
rect 9505 30889 9539 30923
rect 9539 30889 9548 30923
rect 9496 30880 9548 30889
rect 10232 30880 10284 30932
rect 10600 30923 10652 30932
rect 10600 30889 10609 30923
rect 10609 30889 10643 30923
rect 10643 30889 10652 30923
rect 10600 30880 10652 30889
rect 17960 30880 18012 30932
rect 19984 30880 20036 30932
rect 23480 30880 23532 30932
rect 23664 30923 23716 30932
rect 23664 30889 23673 30923
rect 23673 30889 23707 30923
rect 23707 30889 23716 30923
rect 23664 30880 23716 30889
rect 25872 30880 25924 30932
rect 9588 30812 9640 30864
rect 6552 30744 6604 30796
rect 7012 30744 7064 30796
rect 7840 30744 7892 30796
rect 10784 30787 10836 30796
rect 10784 30753 10793 30787
rect 10793 30753 10827 30787
rect 10827 30753 10836 30787
rect 10784 30744 10836 30753
rect 11704 30812 11756 30864
rect 7472 30676 7524 30728
rect 5080 30608 5132 30660
rect 6920 30608 6972 30660
rect 7104 30608 7156 30660
rect 7288 30651 7340 30660
rect 7288 30617 7297 30651
rect 7297 30617 7331 30651
rect 7331 30617 7340 30651
rect 8024 30676 8076 30728
rect 7288 30608 7340 30617
rect 7932 30608 7984 30660
rect 9772 30676 9824 30728
rect 11612 30676 11664 30728
rect 11980 30676 12032 30728
rect 9864 30651 9916 30660
rect 9864 30617 9873 30651
rect 9873 30617 9907 30651
rect 9907 30617 9916 30651
rect 9864 30608 9916 30617
rect 14096 30812 14148 30864
rect 15752 30812 15804 30864
rect 12716 30744 12768 30796
rect 12808 30719 12860 30728
rect 12808 30685 12817 30719
rect 12817 30685 12851 30719
rect 12851 30685 12860 30719
rect 12808 30676 12860 30685
rect 14188 30744 14240 30796
rect 16672 30812 16724 30864
rect 17868 30812 17920 30864
rect 30656 30880 30708 30932
rect 36912 30880 36964 30932
rect 18144 30787 18196 30796
rect 12992 30719 13044 30728
rect 12992 30685 13001 30719
rect 13001 30685 13035 30719
rect 13035 30685 13044 30719
rect 12992 30676 13044 30685
rect 13360 30676 13412 30728
rect 14464 30719 14516 30728
rect 14464 30685 14473 30719
rect 14473 30685 14507 30719
rect 14507 30685 14516 30719
rect 14464 30676 14516 30685
rect 18144 30753 18153 30787
rect 18153 30753 18187 30787
rect 18187 30753 18196 30787
rect 18144 30744 18196 30753
rect 19156 30744 19208 30796
rect 19248 30744 19300 30796
rect 26148 30744 26200 30796
rect 28356 30744 28408 30796
rect 17040 30676 17092 30728
rect 17592 30676 17644 30728
rect 18052 30676 18104 30728
rect 19432 30676 19484 30728
rect 5908 30540 5960 30592
rect 7380 30583 7432 30592
rect 7380 30549 7389 30583
rect 7389 30549 7423 30583
rect 7423 30549 7432 30583
rect 7380 30540 7432 30549
rect 7840 30540 7892 30592
rect 10416 30540 10468 30592
rect 11888 30583 11940 30592
rect 11888 30549 11897 30583
rect 11897 30549 11931 30583
rect 11931 30549 11940 30583
rect 11888 30540 11940 30549
rect 12072 30540 12124 30592
rect 12256 30540 12308 30592
rect 14740 30651 14792 30660
rect 14740 30617 14749 30651
rect 14749 30617 14783 30651
rect 14783 30617 14792 30651
rect 14740 30608 14792 30617
rect 17132 30608 17184 30660
rect 19984 30651 20036 30660
rect 19984 30617 19993 30651
rect 19993 30617 20027 30651
rect 20027 30617 20036 30651
rect 19984 30608 20036 30617
rect 20996 30608 21048 30660
rect 15016 30540 15068 30592
rect 20812 30540 20864 30592
rect 25136 30676 25188 30728
rect 29184 30676 29236 30728
rect 22192 30651 22244 30660
rect 22192 30617 22201 30651
rect 22201 30617 22235 30651
rect 22235 30617 22244 30651
rect 22192 30608 22244 30617
rect 22928 30608 22980 30660
rect 24952 30608 25004 30660
rect 27988 30608 28040 30660
rect 28908 30608 28960 30660
rect 29920 30719 29972 30728
rect 25320 30540 25372 30592
rect 26792 30540 26844 30592
rect 27068 30540 27120 30592
rect 28264 30583 28316 30592
rect 28264 30549 28273 30583
rect 28273 30549 28307 30583
rect 28307 30549 28316 30583
rect 28264 30540 28316 30549
rect 29920 30685 29929 30719
rect 29929 30685 29963 30719
rect 29963 30685 29972 30719
rect 29920 30676 29972 30685
rect 30196 30676 30248 30728
rect 30380 30676 30432 30728
rect 30932 30676 30984 30728
rect 33416 30744 33468 30796
rect 35440 30744 35492 30796
rect 36452 30787 36504 30796
rect 36452 30753 36461 30787
rect 36461 30753 36495 30787
rect 36495 30753 36504 30787
rect 36452 30744 36504 30753
rect 34244 30676 34296 30728
rect 34612 30676 34664 30728
rect 35532 30676 35584 30728
rect 29828 30651 29880 30660
rect 29828 30617 29837 30651
rect 29837 30617 29871 30651
rect 29871 30617 29880 30651
rect 29828 30608 29880 30617
rect 30288 30608 30340 30660
rect 30748 30651 30800 30660
rect 30748 30617 30757 30651
rect 30757 30617 30791 30651
rect 30791 30617 30800 30651
rect 30748 30608 30800 30617
rect 32220 30608 32272 30660
rect 33048 30608 33100 30660
rect 33508 30651 33560 30660
rect 33508 30617 33517 30651
rect 33517 30617 33551 30651
rect 33551 30617 33560 30651
rect 33508 30608 33560 30617
rect 38108 30651 38160 30660
rect 38108 30617 38117 30651
rect 38117 30617 38151 30651
rect 38151 30617 38160 30651
rect 38108 30608 38160 30617
rect 30472 30540 30524 30592
rect 32036 30583 32088 30592
rect 32036 30549 32045 30583
rect 32045 30549 32079 30583
rect 32079 30549 32088 30583
rect 32036 30540 32088 30549
rect 35256 30540 35308 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 6920 30336 6972 30388
rect 8024 30336 8076 30388
rect 10600 30336 10652 30388
rect 12808 30379 12860 30388
rect 12808 30345 12817 30379
rect 12817 30345 12851 30379
rect 12851 30345 12860 30379
rect 12808 30336 12860 30345
rect 14188 30336 14240 30388
rect 14740 30336 14792 30388
rect 7380 30268 7432 30320
rect 12164 30268 12216 30320
rect 13268 30311 13320 30320
rect 5172 30200 5224 30252
rect 5908 30132 5960 30184
rect 7472 30200 7524 30252
rect 7104 30132 7156 30184
rect 4804 30039 4856 30048
rect 4804 30005 4813 30039
rect 4813 30005 4847 30039
rect 4847 30005 4856 30039
rect 4804 29996 4856 30005
rect 4896 29996 4948 30048
rect 7012 30064 7064 30116
rect 8392 30243 8444 30252
rect 8392 30209 8401 30243
rect 8401 30209 8435 30243
rect 8435 30209 8444 30243
rect 8392 30200 8444 30209
rect 9680 30200 9732 30252
rect 9864 30200 9916 30252
rect 10232 30243 10284 30252
rect 10232 30209 10241 30243
rect 10241 30209 10275 30243
rect 10275 30209 10284 30243
rect 10232 30200 10284 30209
rect 11520 30243 11572 30252
rect 11520 30209 11529 30243
rect 11529 30209 11563 30243
rect 11563 30209 11572 30243
rect 11520 30200 11572 30209
rect 11888 30200 11940 30252
rect 12348 30243 12400 30252
rect 12348 30209 12357 30243
rect 12357 30209 12391 30243
rect 12391 30209 12400 30243
rect 12348 30200 12400 30209
rect 13268 30277 13277 30311
rect 13277 30277 13311 30311
rect 13311 30277 13320 30311
rect 13268 30268 13320 30277
rect 13452 30311 13504 30320
rect 13452 30277 13493 30311
rect 13493 30277 13504 30311
rect 15200 30311 15252 30320
rect 13452 30268 13504 30277
rect 15200 30277 15209 30311
rect 15209 30277 15243 30311
rect 15243 30277 15252 30311
rect 15200 30268 15252 30277
rect 15384 30311 15436 30320
rect 15384 30277 15419 30311
rect 15419 30277 15436 30311
rect 15384 30268 15436 30277
rect 14004 30200 14056 30252
rect 14740 30200 14792 30252
rect 15292 30243 15344 30252
rect 10048 30175 10100 30184
rect 10048 30141 10057 30175
rect 10057 30141 10091 30175
rect 10091 30141 10100 30175
rect 10048 30132 10100 30141
rect 11152 30132 11204 30184
rect 8024 30064 8076 30116
rect 11428 30064 11480 30116
rect 11612 30064 11664 30116
rect 12256 30132 12308 30184
rect 12532 30175 12584 30184
rect 12532 30141 12540 30175
rect 12540 30141 12574 30175
rect 12574 30141 12584 30175
rect 15292 30209 15301 30243
rect 15301 30209 15335 30243
rect 15335 30209 15344 30243
rect 15292 30200 15344 30209
rect 19432 30336 19484 30388
rect 19984 30336 20036 30388
rect 16488 30268 16540 30320
rect 17316 30268 17368 30320
rect 20812 30268 20864 30320
rect 20996 30336 21048 30388
rect 22192 30336 22244 30388
rect 22928 30268 22980 30320
rect 27160 30336 27212 30388
rect 29184 30336 29236 30388
rect 30012 30336 30064 30388
rect 30288 30336 30340 30388
rect 27252 30311 27304 30320
rect 27252 30277 27261 30311
rect 27261 30277 27295 30311
rect 27295 30277 27304 30311
rect 27252 30268 27304 30277
rect 27436 30311 27488 30320
rect 27436 30277 27471 30311
rect 27471 30277 27488 30311
rect 27436 30268 27488 30277
rect 27712 30268 27764 30320
rect 29000 30311 29052 30320
rect 29000 30277 29009 30311
rect 29009 30277 29043 30311
rect 29043 30277 29052 30311
rect 29000 30268 29052 30277
rect 18052 30200 18104 30252
rect 18420 30243 18472 30252
rect 18420 30209 18429 30243
rect 18429 30209 18463 30243
rect 18463 30209 18472 30243
rect 18420 30200 18472 30209
rect 18604 30200 18656 30252
rect 19156 30243 19208 30252
rect 19156 30209 19165 30243
rect 19165 30209 19199 30243
rect 19199 30209 19208 30243
rect 19156 30200 19208 30209
rect 19340 30243 19392 30252
rect 19340 30209 19349 30243
rect 19349 30209 19383 30243
rect 19383 30209 19392 30243
rect 19340 30200 19392 30209
rect 12532 30132 12584 30141
rect 15476 30132 15528 30184
rect 15660 30132 15712 30184
rect 16764 30175 16816 30184
rect 16764 30141 16773 30175
rect 16773 30141 16807 30175
rect 16807 30141 16816 30175
rect 16764 30132 16816 30141
rect 18144 30132 18196 30184
rect 18512 30175 18564 30184
rect 18512 30141 18521 30175
rect 18521 30141 18555 30175
rect 18555 30141 18564 30175
rect 18512 30132 18564 30141
rect 19248 30132 19300 30184
rect 19616 30200 19668 30252
rect 20076 30200 20128 30252
rect 20168 30243 20220 30252
rect 20168 30209 20177 30243
rect 20177 30209 20211 30243
rect 20211 30209 20220 30243
rect 20168 30200 20220 30209
rect 20720 30200 20772 30252
rect 22560 30243 22612 30252
rect 22560 30209 22569 30243
rect 22569 30209 22603 30243
rect 22603 30209 22612 30243
rect 22560 30200 22612 30209
rect 23388 30200 23440 30252
rect 24860 30200 24912 30252
rect 28080 30243 28132 30252
rect 22836 30132 22888 30184
rect 24952 30132 25004 30184
rect 26240 30175 26292 30184
rect 26240 30141 26249 30175
rect 26249 30141 26283 30175
rect 26283 30141 26292 30175
rect 26240 30132 26292 30141
rect 18236 30107 18288 30116
rect 9772 29996 9824 30048
rect 11520 29996 11572 30048
rect 11796 29996 11848 30048
rect 11980 29996 12032 30048
rect 13636 30039 13688 30048
rect 13636 30005 13645 30039
rect 13645 30005 13679 30039
rect 13679 30005 13688 30039
rect 13636 29996 13688 30005
rect 13820 29996 13872 30048
rect 18236 30073 18245 30107
rect 18245 30073 18279 30107
rect 18279 30073 18288 30107
rect 18236 30064 18288 30073
rect 17040 29996 17092 30048
rect 17132 29996 17184 30048
rect 26424 30064 26476 30116
rect 28080 30209 28089 30243
rect 28089 30209 28123 30243
rect 28123 30209 28132 30243
rect 28080 30200 28132 30209
rect 30380 30268 30432 30320
rect 30840 30268 30892 30320
rect 31852 30336 31904 30388
rect 32588 30336 32640 30388
rect 35532 30336 35584 30388
rect 31484 30268 31536 30320
rect 35256 30268 35308 30320
rect 37556 30243 37608 30252
rect 27896 30064 27948 30116
rect 29000 30064 29052 30116
rect 19248 29996 19300 30048
rect 26608 29996 26660 30048
rect 27252 29996 27304 30048
rect 27436 29996 27488 30048
rect 27528 29996 27580 30048
rect 37556 30209 37565 30243
rect 37565 30209 37599 30243
rect 37599 30209 37608 30243
rect 37556 30200 37608 30209
rect 30104 30175 30156 30184
rect 30104 30141 30113 30175
rect 30113 30141 30147 30175
rect 30147 30141 30156 30175
rect 30104 30132 30156 30141
rect 34244 30175 34296 30184
rect 29276 30107 29328 30116
rect 29276 30073 29285 30107
rect 29285 30073 29319 30107
rect 29319 30073 29328 30107
rect 29276 30064 29328 30073
rect 31668 30064 31720 30116
rect 32404 30107 32456 30116
rect 32404 30073 32413 30107
rect 32413 30073 32447 30107
rect 32447 30073 32456 30107
rect 32404 30064 32456 30073
rect 32588 30064 32640 30116
rect 34244 30141 34253 30175
rect 34253 30141 34287 30175
rect 34287 30141 34296 30175
rect 34244 30132 34296 30141
rect 33784 30064 33836 30116
rect 31392 29996 31444 30048
rect 31760 29996 31812 30048
rect 34612 29996 34664 30048
rect 36544 30039 36596 30048
rect 36544 30005 36553 30039
rect 36553 30005 36587 30039
rect 36587 30005 36596 30039
rect 36544 29996 36596 30005
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 4896 29792 4948 29844
rect 4804 29588 4856 29640
rect 6184 29631 6236 29640
rect 6184 29597 6193 29631
rect 6193 29597 6227 29631
rect 6227 29597 6236 29631
rect 6184 29588 6236 29597
rect 7012 29588 7064 29640
rect 7472 29656 7524 29708
rect 9128 29656 9180 29708
rect 11060 29656 11112 29708
rect 7564 29631 7616 29640
rect 7564 29597 7573 29631
rect 7573 29597 7607 29631
rect 7607 29597 7616 29631
rect 7564 29588 7616 29597
rect 11336 29631 11388 29640
rect 11336 29597 11345 29631
rect 11345 29597 11379 29631
rect 11379 29597 11388 29631
rect 11336 29588 11388 29597
rect 12808 29792 12860 29844
rect 13452 29792 13504 29844
rect 15752 29792 15804 29844
rect 24860 29792 24912 29844
rect 25412 29792 25464 29844
rect 26792 29835 26844 29844
rect 26792 29801 26801 29835
rect 26801 29801 26835 29835
rect 26835 29801 26844 29835
rect 26792 29792 26844 29801
rect 26976 29835 27028 29844
rect 26976 29801 26985 29835
rect 26985 29801 27019 29835
rect 27019 29801 27028 29835
rect 26976 29792 27028 29801
rect 27988 29835 28040 29844
rect 12348 29767 12400 29776
rect 12348 29733 12357 29767
rect 12357 29733 12391 29767
rect 12391 29733 12400 29767
rect 12348 29724 12400 29733
rect 12624 29724 12676 29776
rect 13636 29724 13688 29776
rect 13452 29656 13504 29708
rect 15108 29656 15160 29708
rect 18328 29699 18380 29708
rect 18328 29665 18337 29699
rect 18337 29665 18371 29699
rect 18371 29665 18380 29699
rect 18328 29656 18380 29665
rect 8024 29520 8076 29572
rect 8576 29520 8628 29572
rect 11428 29563 11480 29572
rect 11428 29529 11437 29563
rect 11437 29529 11471 29563
rect 11471 29529 11480 29563
rect 11428 29520 11480 29529
rect 12072 29520 12124 29572
rect 12256 29520 12308 29572
rect 12624 29631 12676 29640
rect 12624 29597 12633 29631
rect 12633 29597 12667 29631
rect 12667 29597 12676 29631
rect 12624 29588 12676 29597
rect 12992 29588 13044 29640
rect 13636 29588 13688 29640
rect 14740 29631 14792 29640
rect 14740 29597 14749 29631
rect 14749 29597 14783 29631
rect 14783 29597 14792 29631
rect 14740 29588 14792 29597
rect 15016 29588 15068 29640
rect 15660 29588 15712 29640
rect 16396 29588 16448 29640
rect 17224 29588 17276 29640
rect 17960 29631 18012 29640
rect 17960 29597 17969 29631
rect 17969 29597 18003 29631
rect 18003 29597 18012 29631
rect 17960 29588 18012 29597
rect 18144 29631 18196 29640
rect 18144 29597 18150 29631
rect 18150 29597 18196 29631
rect 18144 29588 18196 29597
rect 14188 29520 14240 29572
rect 15384 29520 15436 29572
rect 16120 29520 16172 29572
rect 20168 29656 20220 29708
rect 20812 29699 20864 29708
rect 20812 29665 20821 29699
rect 20821 29665 20855 29699
rect 20855 29665 20864 29699
rect 20812 29656 20864 29665
rect 24400 29656 24452 29708
rect 18696 29588 18748 29640
rect 19340 29588 19392 29640
rect 19616 29631 19668 29640
rect 19616 29597 19625 29631
rect 19625 29597 19659 29631
rect 19659 29597 19668 29631
rect 19616 29588 19668 29597
rect 23388 29588 23440 29640
rect 23664 29631 23716 29640
rect 23664 29597 23673 29631
rect 23673 29597 23707 29631
rect 23707 29597 23716 29631
rect 23664 29588 23716 29597
rect 25412 29588 25464 29640
rect 27712 29724 27764 29776
rect 10232 29452 10284 29504
rect 12440 29452 12492 29504
rect 12900 29452 12952 29504
rect 15936 29452 15988 29504
rect 21088 29563 21140 29572
rect 17316 29495 17368 29504
rect 17316 29461 17325 29495
rect 17325 29461 17359 29495
rect 17359 29461 17368 29495
rect 17316 29452 17368 29461
rect 19156 29452 19208 29504
rect 19248 29452 19300 29504
rect 21088 29529 21097 29563
rect 21097 29529 21131 29563
rect 21131 29529 21140 29563
rect 21088 29520 21140 29529
rect 22652 29520 22704 29572
rect 27344 29588 27396 29640
rect 27620 29631 27672 29640
rect 27620 29597 27629 29631
rect 27629 29597 27663 29631
rect 27663 29597 27672 29631
rect 27620 29588 27672 29597
rect 27988 29801 27997 29835
rect 27997 29801 28031 29835
rect 28031 29801 28040 29835
rect 27988 29792 28040 29801
rect 28264 29792 28316 29844
rect 28172 29724 28224 29776
rect 28908 29792 28960 29844
rect 29276 29792 29328 29844
rect 30104 29835 30156 29844
rect 30104 29801 30113 29835
rect 30113 29801 30147 29835
rect 30147 29801 30156 29835
rect 30104 29792 30156 29801
rect 29920 29724 29972 29776
rect 30288 29724 30340 29776
rect 31024 29724 31076 29776
rect 32036 29792 32088 29844
rect 32956 29792 33008 29844
rect 33508 29792 33560 29844
rect 31484 29699 31536 29708
rect 31484 29665 31493 29699
rect 31493 29665 31527 29699
rect 31527 29665 31536 29699
rect 31484 29656 31536 29665
rect 26056 29520 26108 29572
rect 26608 29563 26660 29572
rect 26608 29529 26617 29563
rect 26617 29529 26651 29563
rect 26651 29529 26660 29563
rect 26608 29520 26660 29529
rect 27528 29520 27580 29572
rect 27896 29520 27948 29572
rect 28816 29563 28868 29572
rect 28816 29529 28825 29563
rect 28825 29529 28859 29563
rect 28859 29529 28868 29563
rect 28816 29520 28868 29529
rect 20996 29452 21048 29504
rect 21824 29452 21876 29504
rect 24768 29452 24820 29504
rect 26700 29452 26752 29504
rect 27988 29452 28040 29504
rect 29092 29452 29144 29504
rect 31668 29588 31720 29640
rect 33232 29631 33284 29640
rect 30656 29520 30708 29572
rect 33232 29597 33241 29631
rect 33241 29597 33275 29631
rect 33275 29597 33284 29631
rect 33232 29588 33284 29597
rect 33416 29631 33468 29640
rect 33416 29597 33425 29631
rect 33425 29597 33459 29631
rect 33459 29597 33468 29631
rect 33416 29588 33468 29597
rect 36084 29656 36136 29708
rect 37464 29656 37516 29708
rect 38108 29699 38160 29708
rect 38108 29665 38117 29699
rect 38117 29665 38151 29699
rect 38151 29665 38160 29699
rect 38108 29656 38160 29665
rect 35532 29631 35584 29640
rect 35532 29597 35541 29631
rect 35541 29597 35575 29631
rect 35575 29597 35584 29631
rect 35532 29588 35584 29597
rect 31392 29452 31444 29504
rect 32128 29452 32180 29504
rect 32312 29452 32364 29504
rect 32588 29495 32640 29504
rect 32588 29461 32615 29495
rect 32615 29461 32640 29495
rect 32588 29452 32640 29461
rect 34704 29563 34756 29572
rect 34704 29529 34713 29563
rect 34713 29529 34747 29563
rect 34747 29529 34756 29563
rect 34704 29520 34756 29529
rect 35348 29520 35400 29572
rect 34520 29452 34572 29504
rect 35900 29452 35952 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 7840 29248 7892 29300
rect 8576 29291 8628 29300
rect 8576 29257 8585 29291
rect 8585 29257 8619 29291
rect 8619 29257 8628 29291
rect 8576 29248 8628 29257
rect 11520 29248 11572 29300
rect 12256 29248 12308 29300
rect 12900 29248 12952 29300
rect 7380 29223 7432 29232
rect 7380 29189 7389 29223
rect 7389 29189 7423 29223
rect 7423 29189 7432 29223
rect 7380 29180 7432 29189
rect 10140 29180 10192 29232
rect 11060 29180 11112 29232
rect 14372 29180 14424 29232
rect 15568 29248 15620 29300
rect 15752 29248 15804 29300
rect 18052 29291 18104 29300
rect 18052 29257 18061 29291
rect 18061 29257 18095 29291
rect 18095 29257 18104 29291
rect 18052 29248 18104 29257
rect 18604 29248 18656 29300
rect 19064 29248 19116 29300
rect 21088 29248 21140 29300
rect 23480 29248 23532 29300
rect 24768 29248 24820 29300
rect 14740 29180 14792 29232
rect 15292 29180 15344 29232
rect 15844 29223 15896 29232
rect 15844 29189 15853 29223
rect 15853 29189 15887 29223
rect 15887 29189 15896 29223
rect 15844 29180 15896 29189
rect 16028 29180 16080 29232
rect 7472 29112 7524 29164
rect 8484 29155 8536 29164
rect 8484 29121 8493 29155
rect 8493 29121 8527 29155
rect 8527 29121 8536 29155
rect 8484 29112 8536 29121
rect 11244 29112 11296 29164
rect 11796 29155 11848 29164
rect 7564 29044 7616 29096
rect 9128 29087 9180 29096
rect 9128 29053 9137 29087
rect 9137 29053 9171 29087
rect 9171 29053 9180 29087
rect 9128 29044 9180 29053
rect 6184 28976 6236 29028
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 12256 29112 12308 29164
rect 12440 29112 12492 29164
rect 12992 29112 13044 29164
rect 13820 29155 13872 29164
rect 11980 29044 12032 29096
rect 13820 29121 13829 29155
rect 13829 29121 13863 29155
rect 13863 29121 13872 29155
rect 13820 29112 13872 29121
rect 14648 29155 14700 29164
rect 14648 29121 14657 29155
rect 14657 29121 14691 29155
rect 14691 29121 14700 29155
rect 14648 29112 14700 29121
rect 15660 29112 15712 29164
rect 16212 29112 16264 29164
rect 16488 29112 16540 29164
rect 15108 29044 15160 29096
rect 17408 29112 17460 29164
rect 18328 29155 18380 29164
rect 18328 29121 18337 29155
rect 18337 29121 18371 29155
rect 18371 29121 18380 29155
rect 18328 29112 18380 29121
rect 23572 29180 23624 29232
rect 24676 29180 24728 29232
rect 25044 29180 25096 29232
rect 25504 29223 25556 29232
rect 25504 29189 25513 29223
rect 25513 29189 25547 29223
rect 25547 29189 25556 29223
rect 25504 29180 25556 29189
rect 19248 29112 19300 29164
rect 20904 29112 20956 29164
rect 21824 29155 21876 29164
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 25596 29112 25648 29164
rect 26056 29112 26108 29164
rect 26976 29112 27028 29164
rect 27160 29248 27212 29300
rect 27712 29248 27764 29300
rect 28448 29248 28500 29300
rect 29920 29248 29972 29300
rect 27252 29223 27304 29232
rect 27252 29189 27261 29223
rect 27261 29189 27295 29223
rect 27295 29189 27304 29223
rect 27252 29180 27304 29189
rect 27160 29155 27212 29164
rect 27160 29121 27169 29155
rect 27169 29121 27203 29155
rect 27203 29121 27212 29155
rect 27160 29112 27212 29121
rect 28540 29155 28592 29164
rect 28540 29121 28549 29155
rect 28549 29121 28583 29155
rect 28583 29121 28592 29155
rect 28540 29112 28592 29121
rect 29184 29180 29236 29232
rect 28816 29112 28868 29164
rect 31024 29248 31076 29300
rect 32220 29248 32272 29300
rect 33232 29180 33284 29232
rect 22008 29087 22060 29096
rect 14924 28976 14976 29028
rect 16120 28976 16172 29028
rect 18512 28976 18564 29028
rect 19524 28976 19576 29028
rect 21180 29019 21232 29028
rect 21180 28985 21189 29019
rect 21189 28985 21223 29019
rect 21223 28985 21232 29019
rect 21180 28976 21232 28985
rect 22008 29053 22017 29087
rect 22017 29053 22051 29087
rect 22051 29053 22060 29087
rect 22008 29044 22060 29053
rect 26516 29044 26568 29096
rect 27620 29044 27672 29096
rect 25136 28976 25188 29028
rect 25964 28976 26016 29028
rect 7472 28908 7524 28960
rect 7748 28951 7800 28960
rect 7748 28917 7757 28951
rect 7757 28917 7791 28951
rect 7791 28917 7800 28951
rect 7748 28908 7800 28917
rect 14372 28908 14424 28960
rect 18420 28908 18472 28960
rect 26240 28908 26292 28960
rect 27068 28976 27120 29028
rect 28724 28976 28776 29028
rect 28908 28976 28960 29028
rect 31392 29155 31444 29164
rect 31392 29121 31401 29155
rect 31401 29121 31435 29155
rect 31435 29121 31444 29155
rect 31392 29112 31444 29121
rect 31760 29112 31812 29164
rect 32128 29155 32180 29164
rect 32128 29121 32137 29155
rect 32137 29121 32171 29155
rect 32171 29121 32180 29155
rect 32128 29112 32180 29121
rect 32312 29155 32364 29164
rect 32312 29121 32321 29155
rect 32321 29121 32355 29155
rect 32355 29121 32364 29155
rect 32312 29112 32364 29121
rect 32956 29155 33008 29164
rect 32956 29121 32965 29155
rect 32965 29121 32999 29155
rect 32999 29121 33008 29155
rect 32956 29112 33008 29121
rect 36544 29180 36596 29232
rect 32864 29044 32916 29096
rect 33140 29087 33192 29096
rect 33140 29053 33149 29087
rect 33149 29053 33183 29087
rect 33183 29053 33192 29087
rect 33140 29044 33192 29053
rect 34244 29112 34296 29164
rect 37556 29155 37608 29164
rect 37556 29121 37565 29155
rect 37565 29121 37599 29155
rect 37599 29121 37608 29155
rect 37556 29112 37608 29121
rect 33692 29044 33744 29096
rect 35348 29044 35400 29096
rect 27252 28908 27304 28960
rect 30564 28908 30616 28960
rect 30932 28908 30984 28960
rect 31484 28908 31536 28960
rect 33784 28908 33836 28960
rect 34060 28908 34112 28960
rect 34152 28908 34204 28960
rect 37924 28908 37976 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 9956 28704 10008 28756
rect 11336 28704 11388 28756
rect 15844 28747 15896 28756
rect 15844 28713 15853 28747
rect 15853 28713 15887 28747
rect 15887 28713 15896 28747
rect 15844 28704 15896 28713
rect 19524 28747 19576 28756
rect 19524 28713 19533 28747
rect 19533 28713 19567 28747
rect 19567 28713 19576 28747
rect 19524 28704 19576 28713
rect 25136 28704 25188 28756
rect 28724 28704 28776 28756
rect 29000 28747 29052 28756
rect 29000 28713 29009 28747
rect 29009 28713 29043 28747
rect 29043 28713 29052 28747
rect 29000 28704 29052 28713
rect 30472 28747 30524 28756
rect 30472 28713 30481 28747
rect 30481 28713 30515 28747
rect 30515 28713 30524 28747
rect 30472 28704 30524 28713
rect 9864 28636 9916 28688
rect 11152 28636 11204 28688
rect 11428 28636 11480 28688
rect 18696 28679 18748 28688
rect 18696 28645 18705 28679
rect 18705 28645 18739 28679
rect 18739 28645 18748 28679
rect 18696 28636 18748 28645
rect 26884 28636 26936 28688
rect 7380 28611 7432 28620
rect 7380 28577 7389 28611
rect 7389 28577 7423 28611
rect 7423 28577 7432 28611
rect 7380 28568 7432 28577
rect 7104 28543 7156 28552
rect 7104 28509 7113 28543
rect 7113 28509 7147 28543
rect 7147 28509 7156 28543
rect 7104 28500 7156 28509
rect 10232 28500 10284 28552
rect 12624 28568 12676 28620
rect 14464 28568 14516 28620
rect 15384 28568 15436 28620
rect 17408 28568 17460 28620
rect 17684 28611 17736 28620
rect 17684 28577 17693 28611
rect 17693 28577 17727 28611
rect 17727 28577 17736 28611
rect 17684 28568 17736 28577
rect 18420 28611 18472 28620
rect 18420 28577 18429 28611
rect 18429 28577 18463 28611
rect 18463 28577 18472 28611
rect 18420 28568 18472 28577
rect 20904 28568 20956 28620
rect 23572 28611 23624 28620
rect 23572 28577 23581 28611
rect 23581 28577 23615 28611
rect 23615 28577 23624 28611
rect 23572 28568 23624 28577
rect 26148 28611 26200 28620
rect 26148 28577 26157 28611
rect 26157 28577 26191 28611
rect 26191 28577 26200 28611
rect 26148 28568 26200 28577
rect 7748 28432 7800 28484
rect 9680 28432 9732 28484
rect 9956 28475 10008 28484
rect 9956 28441 9965 28475
rect 9965 28441 9999 28475
rect 9999 28441 10008 28475
rect 9956 28432 10008 28441
rect 8944 28407 8996 28416
rect 8944 28373 8953 28407
rect 8953 28373 8987 28407
rect 8987 28373 8996 28407
rect 8944 28364 8996 28373
rect 10232 28364 10284 28416
rect 11980 28432 12032 28484
rect 14372 28475 14424 28484
rect 14372 28441 14381 28475
rect 14381 28441 14415 28475
rect 14415 28441 14424 28475
rect 14372 28432 14424 28441
rect 15752 28432 15804 28484
rect 16764 28500 16816 28552
rect 17500 28543 17552 28552
rect 17500 28509 17509 28543
rect 17509 28509 17543 28543
rect 17543 28509 17552 28543
rect 17500 28500 17552 28509
rect 18972 28500 19024 28552
rect 19248 28500 19300 28552
rect 21364 28500 21416 28552
rect 18420 28432 18472 28484
rect 20996 28475 21048 28484
rect 12624 28364 12676 28416
rect 12716 28364 12768 28416
rect 16672 28364 16724 28416
rect 16948 28364 17000 28416
rect 20996 28441 21005 28475
rect 21005 28441 21039 28475
rect 21039 28441 21048 28475
rect 20996 28432 21048 28441
rect 22928 28500 22980 28552
rect 26884 28543 26936 28552
rect 26884 28509 26893 28543
rect 26893 28509 26927 28543
rect 26927 28509 26936 28543
rect 26884 28500 26936 28509
rect 25872 28475 25924 28484
rect 25872 28441 25881 28475
rect 25881 28441 25915 28475
rect 25915 28441 25924 28475
rect 25872 28432 25924 28441
rect 27252 28500 27304 28552
rect 27160 28432 27212 28484
rect 29828 28636 29880 28688
rect 30840 28636 30892 28688
rect 30564 28568 30616 28620
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 29828 28500 29880 28509
rect 30656 28543 30708 28552
rect 30656 28509 30665 28543
rect 30665 28509 30699 28543
rect 30699 28509 30708 28543
rect 30656 28500 30708 28509
rect 30748 28500 30800 28552
rect 31024 28704 31076 28756
rect 31208 28704 31260 28756
rect 31576 28747 31628 28756
rect 31576 28713 31585 28747
rect 31585 28713 31619 28747
rect 31619 28713 31628 28747
rect 31576 28704 31628 28713
rect 31668 28704 31720 28756
rect 33416 28704 33468 28756
rect 34152 28747 34204 28756
rect 34152 28713 34161 28747
rect 34161 28713 34195 28747
rect 34195 28713 34204 28747
rect 34152 28704 34204 28713
rect 34612 28704 34664 28756
rect 33140 28636 33192 28688
rect 31576 28568 31628 28620
rect 31024 28500 31076 28552
rect 32312 28543 32364 28552
rect 32312 28509 32321 28543
rect 32321 28509 32355 28543
rect 32355 28509 32364 28543
rect 32312 28500 32364 28509
rect 33324 28568 33376 28620
rect 34796 28568 34848 28620
rect 35348 28568 35400 28620
rect 37188 28611 37240 28620
rect 37188 28577 37197 28611
rect 37197 28577 37231 28611
rect 37231 28577 37240 28611
rect 37188 28568 37240 28577
rect 37924 28611 37976 28620
rect 37924 28577 37933 28611
rect 37933 28577 37967 28611
rect 37967 28577 37976 28611
rect 37924 28568 37976 28577
rect 33784 28543 33836 28552
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 33784 28500 33836 28509
rect 34520 28500 34572 28552
rect 34980 28500 35032 28552
rect 23572 28364 23624 28416
rect 26332 28364 26384 28416
rect 27528 28364 27580 28416
rect 29000 28364 29052 28416
rect 30196 28364 30248 28416
rect 32496 28407 32548 28416
rect 32496 28373 32505 28407
rect 32505 28373 32539 28407
rect 32539 28373 32548 28407
rect 32496 28364 32548 28373
rect 32680 28475 32732 28484
rect 32680 28441 32689 28475
rect 32689 28441 32723 28475
rect 32723 28441 32732 28475
rect 33692 28475 33744 28484
rect 32680 28432 32732 28441
rect 33692 28441 33709 28475
rect 33709 28441 33744 28475
rect 33692 28432 33744 28441
rect 34060 28432 34112 28484
rect 32772 28364 32824 28416
rect 34796 28364 34848 28416
rect 38108 28543 38160 28552
rect 38108 28509 38117 28543
rect 38117 28509 38151 28543
rect 38151 28509 38160 28543
rect 38108 28500 38160 28509
rect 35716 28364 35768 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 8484 28160 8536 28212
rect 9864 28160 9916 28212
rect 10140 28160 10192 28212
rect 7380 28092 7432 28144
rect 12808 28135 12860 28144
rect 7288 28024 7340 28076
rect 7748 28067 7800 28076
rect 7748 28033 7757 28067
rect 7757 28033 7791 28067
rect 7791 28033 7800 28067
rect 7748 28024 7800 28033
rect 8116 28024 8168 28076
rect 8300 28024 8352 28076
rect 9312 28067 9364 28076
rect 9312 28033 9321 28067
rect 9321 28033 9355 28067
rect 9355 28033 9364 28067
rect 9312 28024 9364 28033
rect 12808 28101 12817 28135
rect 12817 28101 12851 28135
rect 12851 28101 12860 28135
rect 12808 28092 12860 28101
rect 13636 28092 13688 28144
rect 9864 28024 9916 28076
rect 10232 28024 10284 28076
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 9680 27956 9732 28008
rect 11428 27956 11480 28008
rect 6552 27863 6604 27872
rect 6552 27829 6561 27863
rect 6561 27829 6595 27863
rect 6595 27829 6604 27863
rect 6552 27820 6604 27829
rect 7840 27820 7892 27872
rect 9128 27863 9180 27872
rect 9128 27829 9137 27863
rect 9137 27829 9171 27863
rect 9171 27829 9180 27863
rect 9128 27820 9180 27829
rect 12716 28067 12768 28076
rect 12716 28033 12725 28067
rect 12725 28033 12759 28067
rect 12759 28033 12768 28067
rect 12716 28024 12768 28033
rect 12900 28067 12952 28076
rect 12900 28033 12909 28067
rect 12909 28033 12943 28067
rect 12943 28033 12952 28067
rect 12900 28024 12952 28033
rect 13084 28024 13136 28076
rect 13544 28067 13596 28076
rect 13544 28033 13553 28067
rect 13553 28033 13587 28067
rect 13587 28033 13596 28067
rect 13544 28024 13596 28033
rect 12624 27956 12676 28008
rect 14280 28160 14332 28212
rect 14464 28160 14516 28212
rect 15108 28135 15160 28144
rect 15108 28101 15135 28135
rect 15135 28101 15160 28135
rect 15108 28092 15160 28101
rect 15292 28135 15344 28144
rect 15292 28101 15301 28135
rect 15301 28101 15335 28135
rect 15335 28101 15344 28135
rect 15292 28092 15344 28101
rect 15752 28092 15804 28144
rect 17316 28160 17368 28212
rect 17684 28160 17736 28212
rect 20628 28160 20680 28212
rect 21364 28160 21416 28212
rect 22008 28203 22060 28212
rect 22008 28169 22017 28203
rect 22017 28169 22051 28203
rect 22051 28169 22060 28203
rect 22008 28160 22060 28169
rect 22652 28203 22704 28212
rect 22652 28169 22661 28203
rect 22661 28169 22695 28203
rect 22695 28169 22704 28203
rect 22652 28160 22704 28169
rect 25872 28203 25924 28212
rect 25872 28169 25881 28203
rect 25881 28169 25915 28203
rect 25915 28169 25924 28203
rect 25872 28160 25924 28169
rect 16948 28135 17000 28144
rect 16948 28101 16957 28135
rect 16957 28101 16991 28135
rect 16991 28101 17000 28135
rect 16948 28092 17000 28101
rect 18236 28092 18288 28144
rect 22928 28092 22980 28144
rect 27436 28092 27488 28144
rect 27896 28092 27948 28144
rect 14832 28024 14884 28076
rect 15936 28067 15988 28076
rect 15936 28033 15945 28067
rect 15945 28033 15979 28067
rect 15979 28033 15988 28067
rect 15936 28024 15988 28033
rect 16672 28067 16724 28076
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 19248 28067 19300 28076
rect 16948 27956 17000 28008
rect 17500 27956 17552 28008
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 22192 28024 22244 28076
rect 22836 28024 22888 28076
rect 23756 28024 23808 28076
rect 26056 28067 26108 28076
rect 26056 28033 26065 28067
rect 26065 28033 26099 28067
rect 26099 28033 26108 28067
rect 26056 28024 26108 28033
rect 26332 28067 26384 28076
rect 26332 28033 26341 28067
rect 26341 28033 26375 28067
rect 26375 28033 26384 28067
rect 26332 28024 26384 28033
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 27528 28067 27580 28076
rect 9588 27820 9640 27872
rect 12440 27820 12492 27872
rect 12900 27820 12952 27872
rect 13084 27863 13136 27872
rect 13084 27829 13093 27863
rect 13093 27829 13127 27863
rect 13127 27829 13136 27863
rect 13084 27820 13136 27829
rect 14832 27820 14884 27872
rect 14924 27863 14976 27872
rect 14924 27829 14933 27863
rect 14933 27829 14967 27863
rect 14967 27829 14976 27863
rect 14924 27820 14976 27829
rect 15108 27863 15160 27872
rect 15108 27829 15117 27863
rect 15117 27829 15151 27863
rect 15151 27829 15160 27863
rect 19432 27888 19484 27940
rect 18880 27863 18932 27872
rect 15108 27820 15160 27829
rect 18880 27829 18889 27863
rect 18889 27829 18923 27863
rect 18923 27829 18932 27863
rect 18880 27820 18932 27829
rect 21456 27820 21508 27872
rect 21916 27820 21968 27872
rect 23664 27820 23716 27872
rect 24768 27820 24820 27872
rect 25136 27999 25188 28008
rect 25136 27965 25145 27999
rect 25145 27965 25179 27999
rect 25179 27965 25188 27999
rect 26240 27999 26292 28008
rect 25136 27956 25188 27965
rect 26240 27965 26249 27999
rect 26249 27965 26283 27999
rect 26283 27965 26292 27999
rect 27528 28033 27537 28067
rect 27537 28033 27571 28067
rect 27571 28033 27580 28067
rect 27528 28024 27580 28033
rect 26240 27956 26292 27965
rect 25320 27888 25372 27940
rect 26884 27888 26936 27940
rect 30748 28160 30800 28212
rect 29828 28092 29880 28144
rect 29000 28024 29052 28076
rect 30380 28067 30432 28076
rect 30380 28033 30389 28067
rect 30389 28033 30423 28067
rect 30423 28033 30432 28067
rect 30380 28024 30432 28033
rect 32128 28160 32180 28212
rect 32772 28203 32824 28212
rect 32772 28169 32799 28203
rect 32799 28169 32824 28203
rect 32772 28160 32824 28169
rect 32956 28135 33008 28144
rect 32956 28101 32965 28135
rect 32965 28101 32999 28135
rect 32999 28101 33008 28135
rect 32956 28092 33008 28101
rect 33692 28135 33744 28144
rect 31392 28024 31444 28076
rect 31484 28024 31536 28076
rect 33692 28101 33701 28135
rect 33701 28101 33735 28135
rect 33735 28101 33744 28135
rect 33692 28092 33744 28101
rect 34888 28160 34940 28212
rect 34980 28160 35032 28212
rect 33140 28024 33192 28076
rect 33600 28024 33652 28076
rect 29092 27999 29144 28008
rect 29092 27965 29101 27999
rect 29101 27965 29135 27999
rect 29135 27965 29144 27999
rect 29092 27956 29144 27965
rect 30012 27956 30064 28008
rect 31668 27956 31720 28008
rect 33324 27956 33376 28008
rect 28724 27888 28776 27940
rect 30656 27888 30708 27940
rect 31576 27888 31628 27940
rect 32496 27888 32548 27940
rect 30932 27820 30984 27872
rect 31484 27863 31536 27872
rect 31484 27829 31493 27863
rect 31493 27829 31527 27863
rect 31527 27829 31536 27863
rect 31484 27820 31536 27829
rect 33508 27820 33560 27872
rect 35900 28024 35952 28076
rect 38108 28024 38160 28076
rect 34520 27999 34572 28008
rect 34520 27965 34529 27999
rect 34529 27965 34563 27999
rect 34563 27965 34572 27999
rect 34520 27956 34572 27965
rect 34612 27820 34664 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 11704 27616 11756 27668
rect 12808 27616 12860 27668
rect 13084 27616 13136 27668
rect 7012 27548 7064 27600
rect 6184 27480 6236 27532
rect 12256 27548 12308 27600
rect 14464 27548 14516 27600
rect 14924 27548 14976 27600
rect 16764 27616 16816 27668
rect 17408 27616 17460 27668
rect 19248 27659 19300 27668
rect 16856 27548 16908 27600
rect 18144 27548 18196 27600
rect 19248 27625 19257 27659
rect 19257 27625 19291 27659
rect 19291 27625 19300 27659
rect 19248 27616 19300 27625
rect 21916 27616 21968 27668
rect 28172 27616 28224 27668
rect 22284 27548 22336 27600
rect 23756 27591 23808 27600
rect 23756 27557 23765 27591
rect 23765 27557 23799 27591
rect 23799 27557 23808 27591
rect 23756 27548 23808 27557
rect 9588 27523 9640 27532
rect 9588 27489 9597 27523
rect 9597 27489 9631 27523
rect 9631 27489 9640 27523
rect 9588 27480 9640 27489
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 9680 27480 9732 27489
rect 9956 27480 10008 27532
rect 7840 27455 7892 27464
rect 7840 27421 7849 27455
rect 7849 27421 7883 27455
rect 7883 27421 7892 27455
rect 7840 27412 7892 27421
rect 9312 27412 9364 27464
rect 10876 27455 10928 27464
rect 10876 27421 10885 27455
rect 10885 27421 10919 27455
rect 10919 27421 10928 27455
rect 10876 27412 10928 27421
rect 11888 27412 11940 27464
rect 6552 27344 6604 27396
rect 7380 27344 7432 27396
rect 8024 27344 8076 27396
rect 12716 27480 12768 27532
rect 14832 27480 14884 27532
rect 13544 27455 13596 27464
rect 13544 27421 13553 27455
rect 13553 27421 13587 27455
rect 13587 27421 13596 27455
rect 13544 27412 13596 27421
rect 14740 27412 14792 27464
rect 16120 27480 16172 27532
rect 18604 27480 18656 27532
rect 16212 27455 16264 27464
rect 16212 27421 16221 27455
rect 16221 27421 16255 27455
rect 16255 27421 16264 27455
rect 16212 27412 16264 27421
rect 16396 27412 16448 27464
rect 17408 27412 17460 27464
rect 18328 27412 18380 27464
rect 18420 27412 18472 27464
rect 19432 27455 19484 27464
rect 15660 27344 15712 27396
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 7104 27276 7156 27328
rect 9312 27319 9364 27328
rect 9312 27285 9321 27319
rect 9321 27285 9355 27319
rect 9355 27285 9364 27319
rect 9312 27276 9364 27285
rect 14096 27319 14148 27328
rect 14096 27285 14105 27319
rect 14105 27285 14139 27319
rect 14139 27285 14148 27319
rect 14096 27276 14148 27285
rect 16212 27276 16264 27328
rect 18696 27276 18748 27328
rect 19064 27276 19116 27328
rect 20444 27412 20496 27464
rect 20628 27412 20680 27464
rect 23480 27412 23532 27464
rect 23572 27412 23624 27464
rect 27344 27548 27396 27600
rect 27528 27548 27580 27600
rect 28448 27616 28500 27668
rect 31116 27616 31168 27668
rect 31484 27616 31536 27668
rect 32956 27616 33008 27668
rect 28816 27548 28868 27600
rect 24676 27455 24728 27464
rect 24676 27421 24685 27455
rect 24685 27421 24719 27455
rect 24719 27421 24728 27455
rect 24676 27412 24728 27421
rect 25688 27455 25740 27464
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 26056 27412 26108 27464
rect 26332 27455 26384 27464
rect 26332 27421 26341 27455
rect 26341 27421 26375 27455
rect 26375 27421 26384 27455
rect 26332 27412 26384 27421
rect 26792 27412 26844 27464
rect 26976 27412 27028 27464
rect 28080 27480 28132 27532
rect 28172 27480 28224 27532
rect 27528 27455 27580 27464
rect 27528 27421 27537 27455
rect 27537 27421 27571 27455
rect 27571 27421 27580 27455
rect 27528 27412 27580 27421
rect 27712 27412 27764 27464
rect 27804 27412 27856 27464
rect 28448 27455 28500 27464
rect 28448 27421 28457 27455
rect 28457 27421 28491 27455
rect 28491 27421 28500 27455
rect 28448 27412 28500 27421
rect 30748 27548 30800 27600
rect 31116 27480 31168 27532
rect 34612 27548 34664 27600
rect 32680 27480 32732 27532
rect 33508 27480 33560 27532
rect 34428 27480 34480 27532
rect 31208 27455 31260 27464
rect 31208 27421 31217 27455
rect 31217 27421 31251 27455
rect 31251 27421 31260 27455
rect 31208 27412 31260 27421
rect 32588 27455 32640 27464
rect 24584 27344 24636 27396
rect 27436 27387 27488 27396
rect 27436 27353 27445 27387
rect 27445 27353 27479 27387
rect 27479 27353 27488 27387
rect 27436 27344 27488 27353
rect 20352 27276 20404 27328
rect 22744 27319 22796 27328
rect 22744 27285 22753 27319
rect 22753 27285 22787 27319
rect 22787 27285 22796 27319
rect 22744 27276 22796 27285
rect 24676 27276 24728 27328
rect 29736 27344 29788 27396
rect 30380 27344 30432 27396
rect 32588 27421 32597 27455
rect 32597 27421 32631 27455
rect 32631 27421 32640 27455
rect 32588 27412 32640 27421
rect 32956 27412 33008 27464
rect 33600 27344 33652 27396
rect 38660 27480 38712 27532
rect 36268 27455 36320 27464
rect 36268 27421 36277 27455
rect 36277 27421 36311 27455
rect 36311 27421 36320 27455
rect 36268 27412 36320 27421
rect 35532 27344 35584 27396
rect 37372 27344 37424 27396
rect 27896 27276 27948 27328
rect 29092 27276 29144 27328
rect 29552 27276 29604 27328
rect 30564 27276 30616 27328
rect 32128 27276 32180 27328
rect 33508 27276 33560 27328
rect 34704 27276 34756 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9680 27072 9732 27124
rect 11612 27072 11664 27124
rect 11888 27072 11940 27124
rect 14464 27072 14516 27124
rect 14556 27072 14608 27124
rect 18420 27072 18472 27124
rect 18696 27115 18748 27124
rect 18696 27081 18705 27115
rect 18705 27081 18739 27115
rect 18739 27081 18748 27115
rect 18696 27072 18748 27081
rect 18972 27072 19024 27124
rect 7380 27004 7432 27056
rect 9864 27004 9916 27056
rect 6184 26936 6236 26988
rect 11888 26979 11940 26988
rect 11888 26945 11897 26979
rect 11897 26945 11931 26979
rect 11931 26945 11940 26979
rect 11888 26936 11940 26945
rect 6736 26911 6788 26920
rect 6736 26877 6745 26911
rect 6745 26877 6779 26911
rect 6779 26877 6788 26911
rect 6736 26868 6788 26877
rect 8208 26911 8260 26920
rect 8208 26877 8217 26911
rect 8217 26877 8251 26911
rect 8251 26877 8260 26911
rect 8208 26868 8260 26877
rect 9956 26868 10008 26920
rect 10324 26911 10376 26920
rect 10324 26877 10333 26911
rect 10333 26877 10367 26911
rect 10367 26877 10376 26911
rect 10324 26868 10376 26877
rect 13544 27004 13596 27056
rect 14280 27004 14332 27056
rect 14924 27004 14976 27056
rect 15660 26979 15712 26988
rect 9772 26732 9824 26784
rect 14096 26868 14148 26920
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 16212 26936 16264 26988
rect 16948 26979 17000 26988
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 18788 26979 18840 26988
rect 16580 26868 16632 26920
rect 18788 26945 18797 26979
rect 18797 26945 18831 26979
rect 18831 26945 18840 26979
rect 18788 26936 18840 26945
rect 19064 26979 19116 26988
rect 19064 26945 19073 26979
rect 19073 26945 19107 26979
rect 19107 26945 19116 26979
rect 19064 26936 19116 26945
rect 20444 27072 20496 27124
rect 21180 27072 21232 27124
rect 21824 27072 21876 27124
rect 27528 27072 27580 27124
rect 28908 27072 28960 27124
rect 21272 27047 21324 27056
rect 21272 27013 21281 27047
rect 21281 27013 21315 27047
rect 21315 27013 21324 27047
rect 21272 27004 21324 27013
rect 22744 27004 22796 27056
rect 24676 27004 24728 27056
rect 24860 27004 24912 27056
rect 29552 27004 29604 27056
rect 31300 27115 31352 27124
rect 31300 27081 31309 27115
rect 31309 27081 31343 27115
rect 31343 27081 31352 27115
rect 31300 27072 31352 27081
rect 32680 27072 32732 27124
rect 32864 27072 32916 27124
rect 34796 27072 34848 27124
rect 37372 27115 37424 27124
rect 37372 27081 37381 27115
rect 37381 27081 37415 27115
rect 37415 27081 37424 27115
rect 37372 27072 37424 27081
rect 30380 27004 30432 27056
rect 20812 26936 20864 26988
rect 29644 26979 29696 26988
rect 29644 26945 29653 26979
rect 29653 26945 29687 26979
rect 29687 26945 29696 26979
rect 29644 26936 29696 26945
rect 29736 26979 29788 26988
rect 29736 26945 29745 26979
rect 29745 26945 29779 26979
rect 29779 26945 29788 26979
rect 29736 26936 29788 26945
rect 30196 26936 30248 26988
rect 32404 27004 32456 27056
rect 34336 27004 34388 27056
rect 34520 27004 34572 27056
rect 31116 26936 31168 26988
rect 19800 26911 19852 26920
rect 11612 26732 11664 26784
rect 11704 26732 11756 26784
rect 17500 26800 17552 26852
rect 19800 26877 19809 26911
rect 19809 26877 19843 26911
rect 19843 26877 19852 26911
rect 19800 26868 19852 26877
rect 18880 26800 18932 26852
rect 19064 26800 19116 26852
rect 22100 26911 22152 26920
rect 22100 26877 22109 26911
rect 22109 26877 22143 26911
rect 22143 26877 22152 26911
rect 22100 26868 22152 26877
rect 25136 26868 25188 26920
rect 27712 26868 27764 26920
rect 30012 26868 30064 26920
rect 30288 26868 30340 26920
rect 31484 26936 31536 26988
rect 32680 26936 32732 26988
rect 33416 26979 33468 26988
rect 31576 26868 31628 26920
rect 23204 26800 23256 26852
rect 23572 26843 23624 26852
rect 23572 26809 23581 26843
rect 23581 26809 23615 26843
rect 23615 26809 23624 26843
rect 23572 26800 23624 26809
rect 28356 26800 28408 26852
rect 30840 26800 30892 26852
rect 31208 26800 31260 26852
rect 32496 26800 32548 26852
rect 33416 26945 33425 26979
rect 33425 26945 33459 26979
rect 33459 26945 33468 26979
rect 33416 26936 33468 26945
rect 34704 26936 34756 26988
rect 35440 26979 35492 26988
rect 33232 26868 33284 26920
rect 33784 26868 33836 26920
rect 35440 26945 35449 26979
rect 35449 26945 35483 26979
rect 35483 26945 35492 26979
rect 35440 26936 35492 26945
rect 37464 26979 37516 26988
rect 37464 26945 37473 26979
rect 37473 26945 37507 26979
rect 37507 26945 37516 26979
rect 37464 26936 37516 26945
rect 35624 26868 35676 26920
rect 33876 26800 33928 26852
rect 15476 26775 15528 26784
rect 15476 26741 15485 26775
rect 15485 26741 15519 26775
rect 15519 26741 15528 26775
rect 15476 26732 15528 26741
rect 15936 26732 15988 26784
rect 18052 26775 18104 26784
rect 18052 26741 18061 26775
rect 18061 26741 18095 26775
rect 18095 26741 18104 26775
rect 18052 26732 18104 26741
rect 18328 26732 18380 26784
rect 18788 26732 18840 26784
rect 20720 26732 20772 26784
rect 20904 26775 20956 26784
rect 20904 26741 20913 26775
rect 20913 26741 20947 26775
rect 20947 26741 20956 26775
rect 20904 26732 20956 26741
rect 20996 26732 21048 26784
rect 25688 26732 25740 26784
rect 28448 26732 28500 26784
rect 29828 26732 29880 26784
rect 30656 26732 30708 26784
rect 31484 26732 31536 26784
rect 33324 26732 33376 26784
rect 34060 26732 34112 26784
rect 34796 26732 34848 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6736 26528 6788 26580
rect 10324 26528 10376 26580
rect 10876 26528 10928 26580
rect 14556 26528 14608 26580
rect 15384 26528 15436 26580
rect 18052 26528 18104 26580
rect 1860 26324 1912 26376
rect 8208 26435 8260 26444
rect 8208 26401 8217 26435
rect 8217 26401 8251 26435
rect 8251 26401 8260 26435
rect 8208 26392 8260 26401
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 9312 26324 9364 26376
rect 14740 26435 14792 26444
rect 14740 26401 14749 26435
rect 14749 26401 14783 26435
rect 14783 26401 14792 26435
rect 14740 26392 14792 26401
rect 11980 26367 12032 26376
rect 8944 26256 8996 26308
rect 11980 26333 11989 26367
rect 11989 26333 12023 26367
rect 12023 26333 12032 26367
rect 11980 26324 12032 26333
rect 12164 26367 12216 26376
rect 12164 26333 12173 26367
rect 12173 26333 12207 26367
rect 12207 26333 12216 26367
rect 12164 26324 12216 26333
rect 16580 26460 16632 26512
rect 15476 26392 15528 26444
rect 16120 26435 16172 26444
rect 16120 26401 16129 26435
rect 16129 26401 16163 26435
rect 16163 26401 16172 26435
rect 16120 26392 16172 26401
rect 18512 26435 18564 26444
rect 18512 26401 18521 26435
rect 18521 26401 18555 26435
rect 18555 26401 18564 26435
rect 18512 26392 18564 26401
rect 19064 26460 19116 26512
rect 19800 26392 19852 26444
rect 20812 26392 20864 26444
rect 15568 26324 15620 26376
rect 15936 26367 15988 26376
rect 15936 26333 15945 26367
rect 15945 26333 15979 26367
rect 15979 26333 15988 26367
rect 15936 26324 15988 26333
rect 16948 26324 17000 26376
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 18880 26324 18932 26376
rect 21272 26528 21324 26580
rect 24492 26528 24544 26580
rect 25872 26571 25924 26580
rect 25872 26537 25881 26571
rect 25881 26537 25915 26571
rect 25915 26537 25924 26571
rect 25872 26528 25924 26537
rect 26792 26571 26844 26580
rect 26792 26537 26801 26571
rect 26801 26537 26835 26571
rect 26835 26537 26844 26571
rect 26792 26528 26844 26537
rect 22284 26503 22336 26512
rect 22284 26469 22293 26503
rect 22293 26469 22327 26503
rect 22327 26469 22336 26503
rect 22284 26460 22336 26469
rect 27804 26460 27856 26512
rect 28540 26460 28592 26512
rect 25964 26435 26016 26444
rect 25964 26401 25973 26435
rect 25973 26401 26007 26435
rect 26007 26401 26016 26435
rect 25964 26392 26016 26401
rect 21824 26324 21876 26376
rect 22560 26367 22612 26376
rect 22560 26333 22569 26367
rect 22569 26333 22603 26367
rect 22603 26333 22612 26367
rect 22560 26324 22612 26333
rect 12072 26231 12124 26240
rect 12072 26197 12081 26231
rect 12081 26197 12115 26231
rect 12115 26197 12124 26231
rect 12072 26188 12124 26197
rect 15476 26256 15528 26308
rect 15292 26188 15344 26240
rect 17960 26231 18012 26240
rect 17960 26197 17969 26231
rect 17969 26197 18003 26231
rect 18003 26197 18012 26231
rect 17960 26188 18012 26197
rect 20352 26256 20404 26308
rect 21088 26188 21140 26240
rect 22008 26256 22060 26308
rect 24124 26324 24176 26376
rect 24768 26324 24820 26376
rect 26056 26367 26108 26376
rect 26056 26333 26065 26367
rect 26065 26333 26099 26367
rect 26099 26333 26108 26367
rect 26056 26324 26108 26333
rect 23480 26256 23532 26308
rect 24400 26299 24452 26308
rect 24400 26265 24409 26299
rect 24409 26265 24443 26299
rect 24443 26265 24452 26299
rect 24400 26256 24452 26265
rect 25964 26188 26016 26240
rect 28448 26392 28500 26444
rect 28724 26435 28776 26444
rect 28724 26401 28733 26435
rect 28733 26401 28767 26435
rect 28767 26401 28776 26435
rect 28724 26392 28776 26401
rect 29920 26392 29972 26444
rect 26424 26324 26476 26376
rect 26332 26256 26384 26308
rect 27988 26324 28040 26376
rect 27528 26256 27580 26308
rect 27896 26256 27948 26308
rect 28908 26256 28960 26308
rect 30840 26460 30892 26512
rect 32404 26528 32456 26580
rect 34428 26528 34480 26580
rect 30104 26435 30156 26444
rect 30104 26401 30113 26435
rect 30113 26401 30147 26435
rect 30147 26401 30156 26435
rect 30104 26392 30156 26401
rect 30288 26367 30340 26376
rect 30288 26333 30305 26367
rect 30305 26333 30340 26367
rect 30288 26324 30340 26333
rect 30564 26367 30616 26376
rect 30564 26333 30572 26367
rect 30572 26333 30606 26367
rect 30606 26333 30616 26367
rect 30564 26324 30616 26333
rect 31484 26324 31536 26376
rect 32128 26367 32180 26376
rect 32128 26333 32137 26367
rect 32137 26333 32171 26367
rect 32171 26333 32180 26367
rect 32128 26324 32180 26333
rect 34612 26460 34664 26512
rect 33324 26392 33376 26444
rect 33692 26324 33744 26376
rect 34796 26392 34848 26444
rect 33968 26367 34020 26376
rect 33968 26333 33977 26367
rect 33977 26333 34011 26367
rect 34011 26333 34020 26367
rect 33968 26324 34020 26333
rect 34060 26324 34112 26376
rect 30472 26299 30524 26308
rect 30472 26265 30481 26299
rect 30481 26265 30515 26299
rect 30515 26265 30524 26299
rect 32220 26299 32272 26308
rect 30472 26256 30524 26265
rect 32220 26265 32229 26299
rect 32229 26265 32263 26299
rect 32263 26265 32272 26299
rect 32220 26256 32272 26265
rect 32496 26256 32548 26308
rect 33232 26256 33284 26308
rect 33876 26299 33928 26308
rect 33876 26265 33885 26299
rect 33885 26265 33919 26299
rect 33919 26265 33928 26299
rect 35440 26324 35492 26376
rect 35532 26367 35584 26376
rect 35532 26333 35541 26367
rect 35541 26333 35575 26367
rect 35575 26333 35584 26367
rect 35532 26324 35584 26333
rect 35808 26324 35860 26376
rect 36268 26324 36320 26376
rect 37924 26324 37976 26376
rect 35624 26299 35676 26308
rect 33876 26256 33928 26265
rect 35624 26265 35633 26299
rect 35633 26265 35667 26299
rect 35667 26265 35676 26299
rect 35624 26256 35676 26265
rect 30564 26188 30616 26240
rect 30840 26188 30892 26240
rect 37280 26188 37332 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 7380 26027 7432 26036
rect 7380 25993 7389 26027
rect 7389 25993 7423 26027
rect 7423 25993 7432 26027
rect 7380 25984 7432 25993
rect 9864 25984 9916 26036
rect 14280 26027 14332 26036
rect 14280 25993 14289 26027
rect 14289 25993 14323 26027
rect 14323 25993 14332 26027
rect 14280 25984 14332 25993
rect 15568 26027 15620 26036
rect 15568 25993 15577 26027
rect 15577 25993 15611 26027
rect 15611 25993 15620 26027
rect 15568 25984 15620 25993
rect 11796 25916 11848 25968
rect 12072 25916 12124 25968
rect 1860 25891 1912 25900
rect 1860 25857 1869 25891
rect 1869 25857 1903 25891
rect 1903 25857 1912 25891
rect 1860 25848 1912 25857
rect 7288 25891 7340 25900
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 9128 25848 9180 25900
rect 10140 25848 10192 25900
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10232 25848 10284 25857
rect 11612 25848 11664 25900
rect 15292 25916 15344 25968
rect 15476 25916 15528 25968
rect 16396 25916 16448 25968
rect 2780 25780 2832 25832
rect 2872 25823 2924 25832
rect 2872 25789 2881 25823
rect 2881 25789 2915 25823
rect 2915 25789 2924 25823
rect 2872 25780 2924 25789
rect 6552 25780 6604 25832
rect 14832 25848 14884 25900
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 15844 25891 15896 25900
rect 15844 25857 15853 25891
rect 15853 25857 15887 25891
rect 15887 25857 15896 25891
rect 18328 25984 18380 26036
rect 18604 25984 18656 26036
rect 22100 26027 22152 26036
rect 22100 25993 22109 26027
rect 22109 25993 22143 26027
rect 22143 25993 22152 26027
rect 22100 25984 22152 25993
rect 23572 25984 23624 26036
rect 24860 26027 24912 26036
rect 24860 25993 24869 26027
rect 24869 25993 24903 26027
rect 24903 25993 24912 26027
rect 24860 25984 24912 25993
rect 27896 26027 27948 26036
rect 16580 25916 16632 25968
rect 17408 25916 17460 25968
rect 16672 25891 16724 25900
rect 15844 25848 15896 25857
rect 16672 25857 16681 25891
rect 16681 25857 16715 25891
rect 16715 25857 16724 25891
rect 16672 25848 16724 25857
rect 15384 25780 15436 25832
rect 16212 25780 16264 25832
rect 20904 25916 20956 25968
rect 20260 25848 20312 25900
rect 21272 25959 21324 25968
rect 21272 25925 21281 25959
rect 21281 25925 21315 25959
rect 21315 25925 21324 25959
rect 26424 25959 26476 25968
rect 21272 25916 21324 25925
rect 22284 25891 22336 25900
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 22284 25848 22336 25857
rect 22744 25780 22796 25832
rect 20720 25712 20772 25764
rect 20812 25712 20864 25764
rect 21456 25712 21508 25764
rect 23572 25891 23624 25900
rect 23572 25857 23581 25891
rect 23581 25857 23615 25891
rect 23615 25857 23624 25891
rect 24124 25891 24176 25900
rect 23572 25848 23624 25857
rect 24124 25857 24133 25891
rect 24133 25857 24167 25891
rect 24167 25857 24176 25891
rect 24124 25848 24176 25857
rect 24584 25848 24636 25900
rect 25504 25848 25556 25900
rect 26424 25925 26433 25959
rect 26433 25925 26467 25959
rect 26467 25925 26476 25959
rect 26424 25916 26476 25925
rect 26332 25848 26384 25900
rect 25964 25780 26016 25832
rect 26148 25780 26200 25832
rect 27068 25916 27120 25968
rect 27896 25993 27905 26027
rect 27905 25993 27939 26027
rect 27939 25993 27948 26027
rect 27896 25984 27948 25993
rect 30932 25984 30984 26036
rect 31208 25984 31260 26036
rect 32036 25984 32088 26036
rect 33600 25984 33652 26036
rect 33968 25984 34020 26036
rect 35440 25984 35492 26036
rect 30748 25916 30800 25968
rect 31392 25916 31444 25968
rect 34612 25959 34664 25968
rect 34612 25925 34621 25959
rect 34621 25925 34655 25959
rect 34655 25925 34664 25959
rect 34612 25916 34664 25925
rect 35348 25916 35400 25968
rect 28816 25891 28868 25900
rect 28816 25857 28825 25891
rect 28825 25857 28859 25891
rect 28859 25857 28868 25891
rect 28816 25848 28868 25857
rect 29920 25891 29972 25900
rect 29920 25857 29929 25891
rect 29929 25857 29963 25891
rect 29963 25857 29972 25891
rect 29920 25848 29972 25857
rect 30196 25891 30248 25900
rect 30196 25857 30205 25891
rect 30205 25857 30239 25891
rect 30239 25857 30248 25891
rect 30196 25848 30248 25857
rect 30656 25891 30708 25900
rect 30656 25857 30665 25891
rect 30665 25857 30699 25891
rect 30699 25857 30708 25891
rect 30656 25848 30708 25857
rect 31300 25848 31352 25900
rect 31576 25848 31628 25900
rect 32680 25848 32732 25900
rect 34336 25891 34388 25900
rect 23480 25712 23532 25764
rect 25596 25712 25648 25764
rect 28908 25780 28960 25832
rect 30012 25780 30064 25832
rect 30380 25780 30432 25832
rect 30932 25823 30984 25832
rect 30932 25789 30941 25823
rect 30941 25789 30975 25823
rect 30975 25789 30984 25823
rect 30932 25780 30984 25789
rect 32036 25780 32088 25832
rect 33416 25780 33468 25832
rect 34336 25857 34345 25891
rect 34345 25857 34379 25891
rect 34379 25857 34388 25891
rect 34336 25848 34388 25857
rect 37280 25891 37332 25900
rect 37280 25857 37289 25891
rect 37289 25857 37323 25891
rect 37323 25857 37332 25891
rect 37280 25848 37332 25857
rect 37648 25848 37700 25900
rect 35624 25780 35676 25832
rect 28080 25755 28132 25764
rect 28080 25721 28089 25755
rect 28089 25721 28123 25755
rect 28123 25721 28132 25755
rect 28080 25712 28132 25721
rect 9680 25644 9732 25696
rect 13084 25687 13136 25696
rect 13084 25653 13093 25687
rect 13093 25653 13127 25687
rect 13127 25653 13136 25687
rect 13084 25644 13136 25653
rect 18236 25644 18288 25696
rect 19432 25644 19484 25696
rect 20260 25687 20312 25696
rect 20260 25653 20269 25687
rect 20269 25653 20303 25687
rect 20303 25653 20312 25687
rect 20260 25644 20312 25653
rect 20996 25644 21048 25696
rect 22008 25644 22060 25696
rect 25412 25644 25464 25696
rect 26976 25644 27028 25696
rect 27896 25644 27948 25696
rect 36452 25644 36504 25696
rect 38200 25644 38252 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2780 25483 2832 25492
rect 2780 25449 2789 25483
rect 2789 25449 2823 25483
rect 2823 25449 2832 25483
rect 2780 25440 2832 25449
rect 6184 25304 6236 25356
rect 9772 25440 9824 25492
rect 11980 25440 12032 25492
rect 15016 25440 15068 25492
rect 17408 25483 17460 25492
rect 6552 25236 6604 25288
rect 11612 25304 11664 25356
rect 15108 25304 15160 25356
rect 17408 25449 17417 25483
rect 17417 25449 17451 25483
rect 17451 25449 17460 25483
rect 17408 25440 17460 25449
rect 19432 25483 19484 25492
rect 19432 25449 19441 25483
rect 19441 25449 19475 25483
rect 19475 25449 19484 25483
rect 19432 25440 19484 25449
rect 21456 25440 21508 25492
rect 22284 25440 22336 25492
rect 22836 25440 22888 25492
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 20904 25372 20956 25424
rect 23112 25372 23164 25424
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 11060 25236 11112 25288
rect 11888 25236 11940 25288
rect 7564 25168 7616 25220
rect 9864 25211 9916 25220
rect 9864 25177 9898 25211
rect 9898 25177 9916 25211
rect 9864 25168 9916 25177
rect 8208 25100 8260 25152
rect 8484 25100 8536 25152
rect 10140 25100 10192 25152
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 12440 25279 12492 25288
rect 12440 25245 12449 25279
rect 12449 25245 12483 25279
rect 12483 25245 12492 25279
rect 12440 25236 12492 25245
rect 13084 25236 13136 25288
rect 15844 25236 15896 25288
rect 20352 25304 20404 25356
rect 21272 25347 21324 25356
rect 21272 25313 21281 25347
rect 21281 25313 21315 25347
rect 21315 25313 21324 25347
rect 21272 25304 21324 25313
rect 27252 25440 27304 25492
rect 28816 25440 28868 25492
rect 29644 25440 29696 25492
rect 32036 25483 32088 25492
rect 32036 25449 32045 25483
rect 32045 25449 32079 25483
rect 32079 25449 32088 25483
rect 32036 25440 32088 25449
rect 32220 25440 32272 25492
rect 12348 25168 12400 25220
rect 14740 25168 14792 25220
rect 16212 25168 16264 25220
rect 17040 25168 17092 25220
rect 17960 25236 18012 25288
rect 18420 25236 18472 25288
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 20628 25236 20680 25288
rect 20720 25236 20772 25288
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 22744 25279 22796 25288
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 22928 25236 22980 25288
rect 24768 25236 24820 25288
rect 25596 25236 25648 25288
rect 20076 25211 20128 25220
rect 20076 25177 20085 25211
rect 20085 25177 20119 25211
rect 20119 25177 20128 25211
rect 20076 25168 20128 25177
rect 22836 25168 22888 25220
rect 25872 25211 25924 25220
rect 25872 25177 25881 25211
rect 25881 25177 25915 25211
rect 25915 25177 25924 25211
rect 27068 25236 27120 25288
rect 27620 25236 27672 25288
rect 25872 25168 25924 25177
rect 15476 25143 15528 25152
rect 15476 25109 15485 25143
rect 15485 25109 15519 25143
rect 15519 25109 15528 25143
rect 15476 25100 15528 25109
rect 15752 25100 15804 25152
rect 16580 25100 16632 25152
rect 19156 25100 19208 25152
rect 26332 25100 26384 25152
rect 26884 25100 26936 25152
rect 27344 25143 27396 25152
rect 27344 25109 27353 25143
rect 27353 25109 27387 25143
rect 27387 25109 27396 25143
rect 27344 25100 27396 25109
rect 27896 25168 27948 25220
rect 29920 25304 29972 25356
rect 30564 25347 30616 25356
rect 30564 25313 30573 25347
rect 30573 25313 30607 25347
rect 30607 25313 30616 25347
rect 30564 25304 30616 25313
rect 35348 25440 35400 25492
rect 30012 25236 30064 25288
rect 30288 25279 30340 25288
rect 30288 25245 30297 25279
rect 30297 25245 30331 25279
rect 30331 25245 30340 25279
rect 30288 25236 30340 25245
rect 32588 25236 32640 25288
rect 33600 25279 33652 25288
rect 30840 25168 30892 25220
rect 32496 25168 32548 25220
rect 33600 25245 33609 25279
rect 33609 25245 33643 25279
rect 33643 25245 33652 25279
rect 33600 25236 33652 25245
rect 35716 25304 35768 25356
rect 36268 25347 36320 25356
rect 36268 25313 36277 25347
rect 36277 25313 36311 25347
rect 36311 25313 36320 25347
rect 36268 25304 36320 25313
rect 36452 25347 36504 25356
rect 36452 25313 36461 25347
rect 36461 25313 36495 25347
rect 36495 25313 36504 25347
rect 36452 25304 36504 25313
rect 38108 25347 38160 25356
rect 38108 25313 38117 25347
rect 38117 25313 38151 25347
rect 38151 25313 38160 25347
rect 38108 25304 38160 25313
rect 35348 25279 35400 25288
rect 35348 25245 35357 25279
rect 35357 25245 35391 25279
rect 35391 25245 35400 25279
rect 35348 25236 35400 25245
rect 34060 25168 34112 25220
rect 27804 25100 27856 25152
rect 28724 25100 28776 25152
rect 31208 25100 31260 25152
rect 34612 25100 34664 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9128 24896 9180 24948
rect 11796 24896 11848 24948
rect 14740 24939 14792 24948
rect 14740 24905 14749 24939
rect 14749 24905 14783 24939
rect 14783 24905 14792 24939
rect 14740 24896 14792 24905
rect 15476 24896 15528 24948
rect 21272 24896 21324 24948
rect 8300 24871 8352 24880
rect 8300 24837 8309 24871
rect 8309 24837 8343 24871
rect 8343 24837 8352 24871
rect 8300 24828 8352 24837
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7012 24760 7064 24769
rect 9128 24760 9180 24812
rect 10140 24803 10192 24812
rect 7104 24692 7156 24744
rect 9220 24624 9272 24676
rect 10140 24769 10149 24803
rect 10149 24769 10183 24803
rect 10183 24769 10192 24803
rect 10140 24760 10192 24769
rect 12440 24828 12492 24880
rect 12348 24760 12400 24812
rect 13636 24803 13688 24812
rect 12256 24692 12308 24744
rect 13636 24769 13645 24803
rect 13645 24769 13679 24803
rect 13679 24769 13688 24803
rect 13636 24760 13688 24769
rect 13728 24760 13780 24812
rect 16580 24828 16632 24880
rect 19156 24871 19208 24880
rect 19156 24837 19165 24871
rect 19165 24837 19199 24871
rect 19199 24837 19208 24871
rect 19156 24828 19208 24837
rect 20720 24828 20772 24880
rect 24032 24828 24084 24880
rect 27344 24896 27396 24948
rect 28724 24896 28776 24948
rect 30196 24896 30248 24948
rect 30748 24896 30800 24948
rect 31116 24896 31168 24948
rect 28448 24828 28500 24880
rect 14924 24803 14976 24812
rect 14924 24769 14933 24803
rect 14933 24769 14967 24803
rect 14967 24769 14976 24803
rect 14924 24760 14976 24769
rect 17040 24803 17092 24812
rect 11060 24624 11112 24676
rect 11796 24624 11848 24676
rect 17040 24769 17049 24803
rect 17049 24769 17083 24803
rect 17083 24769 17092 24803
rect 17040 24760 17092 24769
rect 21272 24760 21324 24812
rect 21640 24760 21692 24812
rect 21824 24803 21876 24812
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 27160 24803 27212 24812
rect 15568 24692 15620 24744
rect 15752 24735 15804 24744
rect 15752 24701 15761 24735
rect 15761 24701 15795 24735
rect 15795 24701 15804 24735
rect 15752 24692 15804 24701
rect 18512 24692 18564 24744
rect 14464 24624 14516 24676
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 8208 24556 8260 24608
rect 9772 24556 9824 24608
rect 12164 24556 12216 24608
rect 14188 24599 14240 24608
rect 14188 24565 14197 24599
rect 14197 24565 14231 24599
rect 14231 24565 14240 24599
rect 14188 24556 14240 24565
rect 16120 24599 16172 24608
rect 16120 24565 16129 24599
rect 16129 24565 16163 24599
rect 16163 24565 16172 24599
rect 16120 24556 16172 24565
rect 17868 24556 17920 24608
rect 22100 24735 22152 24744
rect 22100 24701 22109 24735
rect 22109 24701 22143 24735
rect 22143 24701 22152 24735
rect 22100 24692 22152 24701
rect 23204 24692 23256 24744
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 25412 24692 25464 24744
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 29736 24760 29788 24812
rect 30656 24828 30708 24880
rect 30380 24803 30432 24812
rect 30380 24769 30389 24803
rect 30389 24769 30423 24803
rect 30423 24769 30432 24803
rect 31576 24828 31628 24880
rect 30380 24760 30432 24769
rect 30932 24803 30984 24812
rect 30932 24769 30941 24803
rect 30941 24769 30975 24803
rect 30975 24769 30984 24803
rect 31116 24803 31168 24812
rect 30932 24760 30984 24769
rect 31116 24769 31125 24803
rect 31125 24769 31159 24803
rect 31159 24769 31168 24803
rect 31116 24760 31168 24769
rect 33508 24760 33560 24812
rect 34336 24803 34388 24812
rect 26148 24735 26200 24744
rect 26148 24701 26157 24735
rect 26157 24701 26191 24735
rect 26191 24701 26200 24735
rect 27712 24735 27764 24744
rect 26148 24692 26200 24701
rect 25964 24624 26016 24676
rect 27712 24701 27721 24735
rect 27721 24701 27755 24735
rect 27755 24701 27764 24735
rect 27712 24692 27764 24701
rect 28356 24692 28408 24744
rect 30288 24692 30340 24744
rect 32404 24735 32456 24744
rect 26700 24624 26752 24676
rect 25136 24556 25188 24608
rect 26148 24556 26200 24608
rect 26424 24556 26476 24608
rect 30472 24624 30524 24676
rect 31392 24556 31444 24608
rect 32036 24556 32088 24608
rect 32404 24701 32413 24735
rect 32413 24701 32447 24735
rect 32447 24701 32456 24735
rect 32404 24692 32456 24701
rect 32956 24692 33008 24744
rect 33784 24692 33836 24744
rect 34336 24769 34345 24803
rect 34345 24769 34379 24803
rect 34379 24769 34388 24803
rect 34336 24760 34388 24769
rect 35716 24760 35768 24812
rect 34612 24735 34664 24744
rect 34336 24624 34388 24676
rect 34612 24701 34621 24735
rect 34621 24701 34655 24735
rect 34655 24701 34664 24735
rect 34612 24692 34664 24701
rect 35808 24692 35860 24744
rect 37280 24624 37332 24676
rect 36268 24556 36320 24608
rect 37832 24599 37884 24608
rect 37832 24565 37841 24599
rect 37841 24565 37875 24599
rect 37875 24565 37884 24599
rect 37832 24556 37884 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 7564 24395 7616 24404
rect 7564 24361 7573 24395
rect 7573 24361 7607 24395
rect 7607 24361 7616 24395
rect 7564 24352 7616 24361
rect 9128 24395 9180 24404
rect 9128 24361 9137 24395
rect 9137 24361 9171 24395
rect 9171 24361 9180 24395
rect 9128 24352 9180 24361
rect 9864 24395 9916 24404
rect 9864 24361 9873 24395
rect 9873 24361 9907 24395
rect 9907 24361 9916 24395
rect 9864 24352 9916 24361
rect 14096 24352 14148 24404
rect 14924 24395 14976 24404
rect 14924 24361 14933 24395
rect 14933 24361 14967 24395
rect 14967 24361 14976 24395
rect 14924 24352 14976 24361
rect 15568 24352 15620 24404
rect 18328 24352 18380 24404
rect 8300 24284 8352 24336
rect 7012 24191 7064 24200
rect 7012 24157 7021 24191
rect 7021 24157 7055 24191
rect 7055 24157 7064 24191
rect 7012 24148 7064 24157
rect 7656 24148 7708 24200
rect 8484 24216 8536 24268
rect 13728 24284 13780 24336
rect 14280 24284 14332 24336
rect 16304 24284 16356 24336
rect 15476 24259 15528 24268
rect 15476 24225 15485 24259
rect 15485 24225 15519 24259
rect 15519 24225 15528 24259
rect 15476 24216 15528 24225
rect 22928 24284 22980 24336
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 9220 24191 9272 24200
rect 9220 24157 9229 24191
rect 9229 24157 9263 24191
rect 9263 24157 9272 24191
rect 9220 24148 9272 24157
rect 9680 24191 9732 24200
rect 9680 24157 9689 24191
rect 9689 24157 9723 24191
rect 9723 24157 9732 24191
rect 9680 24148 9732 24157
rect 9772 24148 9824 24200
rect 11612 24148 11664 24200
rect 12256 24148 12308 24200
rect 7104 24080 7156 24132
rect 6552 24012 6604 24064
rect 9496 24080 9548 24132
rect 11520 24080 11572 24132
rect 12440 24080 12492 24132
rect 16672 24148 16724 24200
rect 17316 24191 17368 24200
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 19248 24191 19300 24200
rect 19248 24157 19257 24191
rect 19257 24157 19291 24191
rect 19291 24157 19300 24191
rect 19248 24148 19300 24157
rect 14372 24123 14424 24132
rect 14372 24089 14381 24123
rect 14381 24089 14415 24123
rect 14415 24089 14424 24123
rect 14372 24080 14424 24089
rect 15752 24080 15804 24132
rect 16120 24080 16172 24132
rect 20168 24080 20220 24132
rect 21180 24216 21232 24268
rect 23572 24352 23624 24404
rect 27160 24352 27212 24404
rect 27896 24395 27948 24404
rect 27896 24361 27905 24395
rect 27905 24361 27939 24395
rect 27939 24361 27948 24395
rect 27896 24352 27948 24361
rect 28356 24395 28408 24404
rect 28356 24361 28365 24395
rect 28365 24361 28399 24395
rect 28399 24361 28408 24395
rect 28356 24352 28408 24361
rect 32496 24395 32548 24404
rect 24032 24284 24084 24336
rect 20628 24080 20680 24132
rect 8484 24012 8536 24064
rect 8576 24012 8628 24064
rect 11888 24012 11940 24064
rect 12164 24012 12216 24064
rect 15568 24012 15620 24064
rect 17776 24012 17828 24064
rect 20996 24012 21048 24064
rect 25780 24216 25832 24268
rect 26424 24259 26476 24268
rect 26424 24225 26433 24259
rect 26433 24225 26467 24259
rect 26467 24225 26476 24259
rect 26424 24216 26476 24225
rect 21824 24191 21876 24200
rect 21824 24157 21833 24191
rect 21833 24157 21867 24191
rect 21867 24157 21876 24191
rect 21824 24148 21876 24157
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 25136 24148 25188 24200
rect 25412 24191 25464 24200
rect 25412 24157 25421 24191
rect 25421 24157 25455 24191
rect 25455 24157 25464 24191
rect 25412 24148 25464 24157
rect 26148 24191 26200 24200
rect 23020 24123 23072 24132
rect 23020 24089 23029 24123
rect 23029 24089 23063 24123
rect 23063 24089 23072 24123
rect 26148 24157 26157 24191
rect 26157 24157 26191 24191
rect 26191 24157 26200 24191
rect 26148 24148 26200 24157
rect 28540 24191 28592 24200
rect 28540 24157 28549 24191
rect 28549 24157 28583 24191
rect 28583 24157 28592 24191
rect 28540 24148 28592 24157
rect 23020 24080 23072 24089
rect 26332 24080 26384 24132
rect 27436 24080 27488 24132
rect 32496 24361 32505 24395
rect 32505 24361 32539 24395
rect 32539 24361 32548 24395
rect 32496 24352 32548 24361
rect 33508 24352 33560 24404
rect 35716 24352 35768 24404
rect 32956 24284 33008 24336
rect 29552 24259 29604 24268
rect 29552 24225 29561 24259
rect 29561 24225 29595 24259
rect 29595 24225 29604 24259
rect 29552 24216 29604 24225
rect 30288 24216 30340 24268
rect 31944 24191 31996 24200
rect 31944 24157 31953 24191
rect 31953 24157 31987 24191
rect 31987 24157 31996 24191
rect 34704 24284 34756 24336
rect 33508 24216 33560 24268
rect 36268 24259 36320 24268
rect 36268 24225 36277 24259
rect 36277 24225 36311 24259
rect 36311 24225 36320 24259
rect 36268 24216 36320 24225
rect 31944 24148 31996 24157
rect 34612 24148 34664 24200
rect 34704 24191 34756 24200
rect 34704 24157 34713 24191
rect 34713 24157 34747 24191
rect 34747 24157 34756 24191
rect 34704 24148 34756 24157
rect 35348 24148 35400 24200
rect 35440 24148 35492 24200
rect 29828 24123 29880 24132
rect 29828 24089 29837 24123
rect 29837 24089 29871 24123
rect 29871 24089 29880 24123
rect 29828 24080 29880 24089
rect 32772 24080 32824 24132
rect 34428 24080 34480 24132
rect 34520 24080 34572 24132
rect 37372 24080 37424 24132
rect 38108 24123 38160 24132
rect 38108 24089 38117 24123
rect 38117 24089 38151 24123
rect 38151 24089 38160 24123
rect 38108 24080 38160 24089
rect 30656 24012 30708 24064
rect 31392 24012 31444 24064
rect 34888 24012 34940 24064
rect 35348 24012 35400 24064
rect 35532 24012 35584 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 6920 23808 6972 23860
rect 7656 23851 7708 23860
rect 7656 23817 7665 23851
rect 7665 23817 7699 23851
rect 7699 23817 7708 23851
rect 7656 23808 7708 23817
rect 7012 23740 7064 23792
rect 7748 23740 7800 23792
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 6644 23715 6696 23724
rect 6644 23681 6653 23715
rect 6653 23681 6687 23715
rect 6687 23681 6696 23715
rect 8300 23808 8352 23860
rect 11520 23851 11572 23860
rect 11520 23817 11529 23851
rect 11529 23817 11563 23851
rect 11563 23817 11572 23851
rect 11520 23808 11572 23817
rect 11888 23808 11940 23860
rect 13360 23808 13412 23860
rect 13636 23808 13688 23860
rect 20076 23808 20128 23860
rect 22100 23808 22152 23860
rect 23756 23808 23808 23860
rect 24124 23851 24176 23860
rect 24124 23817 24133 23851
rect 24133 23817 24167 23851
rect 24167 23817 24176 23851
rect 24124 23808 24176 23817
rect 24676 23808 24728 23860
rect 27252 23808 27304 23860
rect 27436 23808 27488 23860
rect 8208 23740 8260 23792
rect 6644 23672 6696 23681
rect 8852 23715 8904 23724
rect 8852 23681 8861 23715
rect 8861 23681 8895 23715
rect 8895 23681 8904 23715
rect 8852 23672 8904 23681
rect 11612 23740 11664 23792
rect 9680 23672 9732 23724
rect 10140 23672 10192 23724
rect 10416 23715 10468 23724
rect 10416 23681 10425 23715
rect 10425 23681 10459 23715
rect 10459 23681 10468 23715
rect 10416 23672 10468 23681
rect 7104 23604 7156 23656
rect 6736 23536 6788 23588
rect 8484 23604 8536 23656
rect 6368 23511 6420 23520
rect 6368 23477 6377 23511
rect 6377 23477 6411 23511
rect 6411 23477 6420 23511
rect 6368 23468 6420 23477
rect 6920 23468 6972 23520
rect 8116 23468 8168 23520
rect 9404 23511 9456 23520
rect 9404 23477 9413 23511
rect 9413 23477 9447 23511
rect 9447 23477 9456 23511
rect 9404 23468 9456 23477
rect 11796 23681 11805 23708
rect 11805 23681 11839 23708
rect 11839 23681 11848 23708
rect 11796 23656 11848 23681
rect 11980 23715 12032 23724
rect 11980 23681 12015 23715
rect 12015 23681 12032 23715
rect 11980 23672 12032 23681
rect 12164 23715 12216 23724
rect 12164 23681 12173 23715
rect 12173 23681 12207 23715
rect 12207 23681 12216 23715
rect 14648 23740 14700 23792
rect 12164 23672 12216 23681
rect 12900 23672 12952 23724
rect 15292 23715 15344 23724
rect 16580 23740 16632 23792
rect 17224 23740 17276 23792
rect 17316 23740 17368 23792
rect 17868 23740 17920 23792
rect 15292 23681 15320 23715
rect 15320 23681 15344 23715
rect 15292 23672 15344 23681
rect 16672 23715 16724 23724
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 11888 23536 11940 23588
rect 10600 23468 10652 23520
rect 19248 23672 19300 23724
rect 19984 23672 20036 23724
rect 20536 23715 20588 23724
rect 20536 23681 20545 23715
rect 20545 23681 20579 23715
rect 20579 23681 20588 23715
rect 20536 23672 20588 23681
rect 20628 23672 20680 23724
rect 23388 23672 23440 23724
rect 23848 23672 23900 23724
rect 24584 23715 24636 23724
rect 20352 23604 20404 23656
rect 22100 23647 22152 23656
rect 22100 23613 22109 23647
rect 22109 23613 22143 23647
rect 22143 23613 22152 23647
rect 22100 23604 22152 23613
rect 23664 23604 23716 23656
rect 24584 23681 24593 23715
rect 24593 23681 24627 23715
rect 24627 23681 24636 23715
rect 24584 23672 24636 23681
rect 24676 23672 24728 23724
rect 26332 23740 26384 23792
rect 25596 23647 25648 23656
rect 25596 23613 25605 23647
rect 25605 23613 25639 23647
rect 25639 23613 25648 23647
rect 25596 23604 25648 23613
rect 12072 23536 12124 23588
rect 12532 23536 12584 23588
rect 14096 23536 14148 23588
rect 31024 23672 31076 23724
rect 32772 23808 32824 23860
rect 34520 23808 34572 23860
rect 34888 23808 34940 23860
rect 37372 23851 37424 23860
rect 33508 23715 33560 23724
rect 33508 23681 33517 23715
rect 33517 23681 33551 23715
rect 33551 23681 33560 23715
rect 33508 23672 33560 23681
rect 34336 23740 34388 23792
rect 37372 23817 37381 23851
rect 37381 23817 37415 23851
rect 37415 23817 37424 23851
rect 37372 23808 37424 23817
rect 35348 23672 35400 23724
rect 37280 23715 37332 23724
rect 13176 23468 13228 23520
rect 17500 23468 17552 23520
rect 20168 23468 20220 23520
rect 23296 23468 23348 23520
rect 23756 23468 23808 23520
rect 33692 23604 33744 23656
rect 34336 23604 34388 23656
rect 37280 23681 37289 23715
rect 37289 23681 37323 23715
rect 37323 23681 37332 23715
rect 37280 23672 37332 23681
rect 37464 23604 37516 23656
rect 31944 23536 31996 23588
rect 36084 23536 36136 23588
rect 35716 23511 35768 23520
rect 35716 23477 35725 23511
rect 35725 23477 35759 23511
rect 35759 23477 35768 23511
rect 35716 23468 35768 23477
rect 36360 23511 36412 23520
rect 36360 23477 36369 23511
rect 36369 23477 36403 23511
rect 36403 23477 36412 23511
rect 36360 23468 36412 23477
rect 36544 23468 36596 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8852 23264 8904 23316
rect 7748 23171 7800 23180
rect 7748 23137 7757 23171
rect 7757 23137 7791 23171
rect 7791 23137 7800 23171
rect 7748 23128 7800 23137
rect 10416 23264 10468 23316
rect 12348 23264 12400 23316
rect 12900 23307 12952 23316
rect 12900 23273 12909 23307
rect 12909 23273 12943 23307
rect 12943 23273 12952 23307
rect 12900 23264 12952 23273
rect 4344 23060 4396 23112
rect 4620 23060 4672 23112
rect 6368 23060 6420 23112
rect 7840 23060 7892 23112
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 10416 23060 10468 23112
rect 11980 23128 12032 23180
rect 8760 22992 8812 23044
rect 12348 23060 12400 23112
rect 14188 23128 14240 23180
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 13360 23103 13412 23112
rect 13360 23069 13395 23103
rect 13395 23069 13412 23103
rect 13360 23060 13412 23069
rect 13820 23060 13872 23112
rect 14096 23060 14148 23112
rect 16856 23307 16908 23316
rect 16856 23273 16865 23307
rect 16865 23273 16899 23307
rect 16899 23273 16908 23307
rect 16856 23264 16908 23273
rect 19064 23264 19116 23316
rect 21456 23307 21508 23316
rect 21456 23273 21465 23307
rect 21465 23273 21499 23307
rect 21499 23273 21508 23307
rect 21456 23264 21508 23273
rect 22100 23264 22152 23316
rect 34520 23264 34572 23316
rect 35440 23307 35492 23316
rect 35440 23273 35449 23307
rect 35449 23273 35483 23307
rect 35483 23273 35492 23307
rect 35440 23264 35492 23273
rect 17040 23196 17092 23248
rect 19432 23196 19484 23248
rect 15476 23128 15528 23180
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 11888 23035 11940 23044
rect 11888 23001 11897 23035
rect 11897 23001 11931 23035
rect 11931 23001 11940 23035
rect 11888 22992 11940 23001
rect 13176 23035 13228 23044
rect 13176 23001 13185 23035
rect 13185 23001 13219 23035
rect 13219 23001 13228 23035
rect 13176 22992 13228 23001
rect 10784 22924 10836 22976
rect 11428 22967 11480 22976
rect 11428 22933 11437 22967
rect 11437 22933 11471 22967
rect 11471 22933 11480 22967
rect 11428 22924 11480 22933
rect 12164 22924 12216 22976
rect 14004 22992 14056 23044
rect 15476 23035 15528 23044
rect 15476 23001 15485 23035
rect 15485 23001 15519 23035
rect 15519 23001 15528 23035
rect 15476 22992 15528 23001
rect 14556 22924 14608 22976
rect 16396 23128 16448 23180
rect 15752 23103 15804 23112
rect 15752 23069 15761 23103
rect 15761 23069 15795 23103
rect 15795 23069 15804 23103
rect 15752 23060 15804 23069
rect 16764 23060 16816 23112
rect 17040 23060 17092 23112
rect 20536 23128 20588 23180
rect 24584 23196 24636 23248
rect 25596 23196 25648 23248
rect 23388 23128 23440 23180
rect 17500 23103 17552 23112
rect 17500 23069 17509 23103
rect 17509 23069 17543 23103
rect 17543 23069 17552 23103
rect 17960 23103 18012 23112
rect 17500 23060 17552 23069
rect 17960 23069 17969 23103
rect 17969 23069 18003 23103
rect 18003 23069 18012 23103
rect 17960 23060 18012 23069
rect 18236 23060 18288 23112
rect 19432 23060 19484 23112
rect 20076 23060 20128 23112
rect 20168 23060 20220 23112
rect 21180 23103 21232 23112
rect 21180 23069 21189 23103
rect 21189 23069 21223 23103
rect 21223 23069 21232 23103
rect 21180 23060 21232 23069
rect 21364 23060 21416 23112
rect 26240 23128 26292 23180
rect 29552 23171 29604 23180
rect 25044 23060 25096 23112
rect 25412 23060 25464 23112
rect 27068 23103 27120 23112
rect 27068 23069 27077 23103
rect 27077 23069 27111 23103
rect 27111 23069 27120 23103
rect 27068 23060 27120 23069
rect 29552 23137 29561 23171
rect 29561 23137 29595 23171
rect 29595 23137 29604 23171
rect 29552 23128 29604 23137
rect 30840 23196 30892 23248
rect 32036 23171 32088 23180
rect 23388 22992 23440 23044
rect 24584 23035 24636 23044
rect 24584 23001 24593 23035
rect 24593 23001 24627 23035
rect 24627 23001 24636 23035
rect 24584 22992 24636 23001
rect 24952 23035 25004 23044
rect 24952 23001 24961 23035
rect 24961 23001 24995 23035
rect 24995 23001 25004 23035
rect 24952 22992 25004 23001
rect 15660 22924 15712 22976
rect 17224 22924 17276 22976
rect 18052 22967 18104 22976
rect 18052 22933 18061 22967
rect 18061 22933 18095 22967
rect 18095 22933 18104 22967
rect 18052 22924 18104 22933
rect 18880 22924 18932 22976
rect 20444 22924 20496 22976
rect 24308 22924 24360 22976
rect 24492 22924 24544 22976
rect 25780 22992 25832 23044
rect 29460 22992 29512 23044
rect 30380 22992 30432 23044
rect 32036 23137 32045 23171
rect 32045 23137 32079 23171
rect 32079 23137 32088 23171
rect 32036 23128 32088 23137
rect 36360 23171 36412 23180
rect 33416 23060 33468 23112
rect 36360 23137 36369 23171
rect 36369 23137 36403 23171
rect 36403 23137 36412 23171
rect 36360 23128 36412 23137
rect 38016 23171 38068 23180
rect 38016 23137 38025 23171
rect 38025 23137 38059 23171
rect 38059 23137 38068 23171
rect 38016 23128 38068 23137
rect 31852 22992 31904 23044
rect 32312 23035 32364 23044
rect 32312 23001 32321 23035
rect 32321 23001 32355 23035
rect 32355 23001 32364 23035
rect 32312 22992 32364 23001
rect 25504 22967 25556 22976
rect 25504 22933 25513 22967
rect 25513 22933 25547 22967
rect 25547 22933 25556 22967
rect 25504 22924 25556 22933
rect 26516 22967 26568 22976
rect 26516 22933 26525 22967
rect 26525 22933 26559 22967
rect 26559 22933 26568 22967
rect 26516 22924 26568 22933
rect 27252 22967 27304 22976
rect 27252 22933 27261 22967
rect 27261 22933 27295 22967
rect 27295 22933 27304 22967
rect 27252 22924 27304 22933
rect 27804 22967 27856 22976
rect 27804 22933 27813 22967
rect 27813 22933 27847 22967
rect 27847 22933 27856 22967
rect 27804 22924 27856 22933
rect 31300 22967 31352 22976
rect 31300 22933 31309 22967
rect 31309 22933 31343 22967
rect 31343 22933 31352 22967
rect 31300 22924 31352 22933
rect 33048 22924 33100 22976
rect 35992 23060 36044 23112
rect 36176 22924 36228 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 8760 22763 8812 22772
rect 8760 22729 8769 22763
rect 8769 22729 8803 22763
rect 8803 22729 8812 22763
rect 8760 22720 8812 22729
rect 9404 22720 9456 22772
rect 9680 22720 9732 22772
rect 7840 22652 7892 22704
rect 11980 22720 12032 22772
rect 12256 22720 12308 22772
rect 12532 22763 12584 22772
rect 12532 22729 12541 22763
rect 12541 22729 12575 22763
rect 12575 22729 12584 22763
rect 12532 22720 12584 22729
rect 13176 22720 13228 22772
rect 16948 22720 17000 22772
rect 24308 22720 24360 22772
rect 29460 22763 29512 22772
rect 11428 22652 11480 22704
rect 4344 22627 4396 22636
rect 4344 22593 4353 22627
rect 4353 22593 4387 22627
rect 4387 22593 4396 22627
rect 4344 22584 4396 22593
rect 6552 22627 6604 22636
rect 6552 22593 6561 22627
rect 6561 22593 6595 22627
rect 6595 22593 6604 22627
rect 6552 22584 6604 22593
rect 6644 22627 6696 22636
rect 6644 22593 6653 22627
rect 6653 22593 6687 22627
rect 6687 22593 6696 22627
rect 6644 22584 6696 22593
rect 6828 22627 6880 22636
rect 6828 22593 6863 22627
rect 6863 22593 6880 22627
rect 6828 22584 6880 22593
rect 7012 22559 7064 22568
rect 7012 22525 7021 22559
rect 7021 22525 7055 22559
rect 7055 22525 7064 22559
rect 7012 22516 7064 22525
rect 7748 22584 7800 22636
rect 8300 22584 8352 22636
rect 8392 22516 8444 22568
rect 8576 22627 8628 22636
rect 8576 22593 8585 22627
rect 8585 22593 8619 22627
rect 8619 22593 8628 22627
rect 8576 22584 8628 22593
rect 7564 22448 7616 22500
rect 8484 22448 8536 22500
rect 10140 22584 10192 22636
rect 10784 22627 10836 22636
rect 10784 22593 10793 22627
rect 10793 22593 10827 22627
rect 10827 22593 10836 22627
rect 10784 22584 10836 22593
rect 11244 22516 11296 22568
rect 12164 22584 12216 22636
rect 12716 22559 12768 22568
rect 5908 22380 5960 22432
rect 8300 22423 8352 22432
rect 8300 22389 8309 22423
rect 8309 22389 8343 22423
rect 8343 22389 8352 22423
rect 8300 22380 8352 22389
rect 8852 22380 8904 22432
rect 10416 22448 10468 22500
rect 11152 22448 11204 22500
rect 12716 22525 12725 22559
rect 12725 22525 12759 22559
rect 12759 22525 12768 22559
rect 12716 22516 12768 22525
rect 13636 22652 13688 22704
rect 14464 22695 14516 22704
rect 14464 22661 14473 22695
rect 14473 22661 14507 22695
rect 14507 22661 14516 22695
rect 14464 22652 14516 22661
rect 15752 22652 15804 22704
rect 16212 22652 16264 22704
rect 13820 22584 13872 22636
rect 14004 22627 14056 22636
rect 14004 22593 14013 22627
rect 14013 22593 14047 22627
rect 14047 22593 14056 22627
rect 14004 22584 14056 22593
rect 14372 22584 14424 22636
rect 15660 22627 15712 22636
rect 15660 22593 15669 22627
rect 15669 22593 15703 22627
rect 15703 22593 15712 22627
rect 15660 22584 15712 22593
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 16120 22584 16172 22593
rect 17500 22652 17552 22704
rect 18880 22695 18932 22704
rect 18880 22661 18889 22695
rect 18889 22661 18923 22695
rect 18923 22661 18932 22695
rect 18880 22652 18932 22661
rect 19892 22652 19944 22704
rect 17224 22627 17276 22636
rect 17224 22593 17233 22627
rect 17233 22593 17267 22627
rect 17267 22593 17276 22627
rect 17224 22584 17276 22593
rect 18144 22627 18196 22636
rect 18144 22593 18153 22627
rect 18153 22593 18187 22627
rect 18187 22593 18196 22627
rect 18144 22584 18196 22593
rect 22744 22652 22796 22704
rect 25504 22652 25556 22704
rect 21364 22584 21416 22636
rect 29460 22729 29469 22763
rect 29469 22729 29503 22763
rect 29503 22729 29512 22763
rect 29460 22720 29512 22729
rect 33416 22720 33468 22772
rect 27252 22695 27304 22704
rect 27252 22661 27261 22695
rect 27261 22661 27295 22695
rect 27295 22661 27304 22695
rect 27252 22652 27304 22661
rect 27804 22652 27856 22704
rect 10692 22423 10744 22432
rect 10692 22389 10701 22423
rect 10701 22389 10735 22423
rect 10735 22389 10744 22423
rect 10692 22380 10744 22389
rect 12348 22380 12400 22432
rect 19432 22516 19484 22568
rect 19984 22559 20036 22568
rect 19984 22525 19993 22559
rect 19993 22525 20027 22559
rect 20027 22525 20036 22559
rect 19984 22516 20036 22525
rect 22284 22516 22336 22568
rect 16672 22448 16724 22500
rect 22560 22448 22612 22500
rect 22652 22448 22704 22500
rect 23204 22516 23256 22568
rect 23572 22516 23624 22568
rect 23664 22448 23716 22500
rect 15292 22380 15344 22432
rect 19340 22380 19392 22432
rect 19616 22423 19668 22432
rect 19616 22389 19625 22423
rect 19625 22389 19659 22423
rect 19659 22389 19668 22423
rect 19616 22380 19668 22389
rect 21180 22380 21232 22432
rect 23020 22380 23072 22432
rect 25504 22423 25556 22432
rect 25504 22389 25513 22423
rect 25513 22389 25547 22423
rect 25547 22389 25556 22423
rect 25504 22380 25556 22389
rect 26148 22448 26200 22500
rect 29276 22627 29328 22636
rect 29276 22593 29285 22627
rect 29285 22593 29319 22627
rect 29319 22593 29328 22627
rect 29276 22584 29328 22593
rect 30104 22627 30156 22636
rect 30104 22593 30113 22627
rect 30113 22593 30147 22627
rect 30147 22593 30156 22627
rect 30104 22584 30156 22593
rect 30472 22584 30524 22636
rect 30840 22584 30892 22636
rect 29000 22380 29052 22432
rect 30012 22423 30064 22432
rect 30012 22389 30021 22423
rect 30021 22389 30055 22423
rect 30055 22389 30064 22423
rect 30012 22380 30064 22389
rect 30104 22380 30156 22432
rect 33876 22516 33928 22568
rect 31944 22448 31996 22500
rect 33784 22448 33836 22500
rect 34612 22584 34664 22636
rect 37464 22584 37516 22636
rect 36544 22516 36596 22568
rect 36728 22559 36780 22568
rect 36728 22525 36737 22559
rect 36737 22525 36771 22559
rect 36771 22525 36780 22559
rect 36728 22516 36780 22525
rect 37004 22516 37056 22568
rect 32128 22380 32180 22432
rect 34704 22380 34756 22432
rect 36452 22448 36504 22500
rect 37280 22380 37332 22432
rect 37924 22380 37976 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 7104 22176 7156 22228
rect 7656 22108 7708 22160
rect 8300 22176 8352 22228
rect 10416 22219 10468 22228
rect 10416 22185 10425 22219
rect 10425 22185 10459 22219
rect 10459 22185 10468 22219
rect 10416 22176 10468 22185
rect 10600 22176 10652 22228
rect 10692 22176 10744 22228
rect 14188 22176 14240 22228
rect 14648 22176 14700 22228
rect 17960 22176 18012 22228
rect 20536 22176 20588 22228
rect 25044 22219 25096 22228
rect 25044 22185 25053 22219
rect 25053 22185 25087 22219
rect 25087 22185 25096 22219
rect 25044 22176 25096 22185
rect 33048 22219 33100 22228
rect 5908 22040 5960 22092
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 6736 21972 6788 22024
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 11336 22108 11388 22160
rect 11980 22108 12032 22160
rect 10692 22040 10744 22092
rect 7012 21972 7064 21981
rect 8116 21972 8168 22024
rect 10232 21972 10284 22024
rect 10784 21972 10836 22024
rect 11244 21972 11296 22024
rect 11336 22015 11388 22024
rect 11336 21981 11345 22015
rect 11345 21981 11379 22015
rect 11379 21981 11388 22015
rect 11520 22015 11572 22024
rect 11336 21972 11388 21981
rect 11520 21981 11529 22015
rect 11529 21981 11563 22015
rect 11563 21981 11572 22015
rect 11520 21972 11572 21981
rect 11888 22040 11940 22092
rect 14464 22108 14516 22160
rect 16396 22108 16448 22160
rect 13084 22040 13136 22092
rect 15752 22083 15804 22092
rect 15752 22049 15761 22083
rect 15761 22049 15795 22083
rect 15795 22049 15804 22083
rect 15752 22040 15804 22049
rect 12348 21972 12400 22024
rect 13636 21972 13688 22024
rect 15476 21972 15528 22024
rect 7748 21879 7800 21888
rect 7748 21845 7757 21879
rect 7757 21845 7791 21879
rect 7791 21845 7800 21879
rect 7748 21836 7800 21845
rect 8760 21904 8812 21956
rect 15844 21904 15896 21956
rect 16672 22015 16724 22024
rect 16672 21981 16681 22015
rect 16681 21981 16715 22015
rect 16715 21981 16724 22015
rect 18236 22040 18288 22092
rect 16672 21972 16724 21981
rect 17132 21972 17184 22024
rect 19156 21972 19208 22024
rect 19616 22108 19668 22160
rect 23572 22108 23624 22160
rect 19892 22083 19944 22092
rect 19892 22049 19901 22083
rect 19901 22049 19935 22083
rect 19935 22049 19944 22083
rect 19892 22040 19944 22049
rect 21364 22040 21416 22092
rect 22284 22015 22336 22024
rect 16396 21904 16448 21956
rect 18420 21947 18472 21956
rect 18420 21913 18429 21947
rect 18429 21913 18463 21947
rect 18463 21913 18472 21947
rect 18420 21904 18472 21913
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 22744 21947 22796 21956
rect 22744 21913 22753 21947
rect 22753 21913 22787 21947
rect 22787 21913 22796 21947
rect 22744 21904 22796 21913
rect 23020 21904 23072 21956
rect 26148 22040 26200 22092
rect 27712 22040 27764 22092
rect 29552 22108 29604 22160
rect 33048 22185 33057 22219
rect 33057 22185 33091 22219
rect 33091 22185 33100 22219
rect 33048 22176 33100 22185
rect 33784 22219 33836 22228
rect 33784 22185 33793 22219
rect 33793 22185 33827 22219
rect 33827 22185 33836 22219
rect 33784 22176 33836 22185
rect 35716 22176 35768 22228
rect 35992 22176 36044 22228
rect 37188 22176 37240 22228
rect 35440 22108 35492 22160
rect 23296 21972 23348 22024
rect 23664 21972 23716 22024
rect 25504 21972 25556 22024
rect 27988 21972 28040 22024
rect 31116 22040 31168 22092
rect 28356 22015 28408 22024
rect 28356 21981 28365 22015
rect 28365 21981 28399 22015
rect 28399 21981 28408 22015
rect 28356 21972 28408 21981
rect 29092 21972 29144 22024
rect 30104 21972 30156 22024
rect 35900 22040 35952 22092
rect 37464 22083 37516 22092
rect 37464 22049 37473 22083
rect 37473 22049 37507 22083
rect 37507 22049 37516 22083
rect 37464 22040 37516 22049
rect 37924 22083 37976 22092
rect 37924 22049 37933 22083
rect 37933 22049 37967 22083
rect 37967 22049 37976 22083
rect 37924 22040 37976 22049
rect 38200 22040 38252 22092
rect 34796 21972 34848 22024
rect 24952 21904 25004 21956
rect 26332 21904 26384 21956
rect 26516 21904 26568 21956
rect 30380 21904 30432 21956
rect 30748 21947 30800 21956
rect 30748 21913 30757 21947
rect 30757 21913 30791 21947
rect 30791 21913 30800 21947
rect 30748 21904 30800 21913
rect 32128 21904 32180 21956
rect 35348 21947 35400 21956
rect 11612 21836 11664 21888
rect 14832 21836 14884 21888
rect 19248 21879 19300 21888
rect 19248 21845 19257 21879
rect 19257 21845 19291 21879
rect 19291 21845 19300 21879
rect 19248 21836 19300 21845
rect 19432 21836 19484 21888
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20076 21836 20128 21845
rect 23848 21836 23900 21888
rect 24400 21879 24452 21888
rect 24400 21845 24409 21879
rect 24409 21845 24443 21879
rect 24443 21845 24452 21879
rect 24400 21836 24452 21845
rect 24584 21836 24636 21888
rect 26240 21836 26292 21888
rect 27620 21836 27672 21888
rect 28908 21879 28960 21888
rect 28908 21845 28917 21879
rect 28917 21845 28951 21879
rect 28951 21845 28960 21879
rect 28908 21836 28960 21845
rect 32220 21879 32272 21888
rect 32220 21845 32229 21879
rect 32229 21845 32263 21879
rect 32263 21845 32272 21879
rect 35348 21913 35357 21947
rect 35357 21913 35391 21947
rect 35391 21913 35400 21947
rect 35348 21904 35400 21913
rect 37280 21904 37332 21956
rect 33232 21879 33284 21888
rect 32220 21836 32272 21845
rect 33232 21845 33241 21879
rect 33241 21845 33275 21879
rect 33275 21845 33284 21879
rect 33232 21836 33284 21845
rect 33968 21879 34020 21888
rect 33968 21845 33995 21879
rect 33995 21845 34020 21879
rect 33968 21836 34020 21845
rect 34060 21836 34112 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4620 21632 4672 21684
rect 6368 21632 6420 21684
rect 7564 21632 7616 21684
rect 8024 21607 8076 21616
rect 8024 21573 8033 21607
rect 8033 21573 8067 21607
rect 8067 21573 8076 21607
rect 8024 21564 8076 21573
rect 8392 21564 8444 21616
rect 6368 21539 6420 21548
rect 6368 21505 6377 21539
rect 6377 21505 6411 21539
rect 6411 21505 6420 21539
rect 6368 21496 6420 21505
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 6644 21471 6696 21480
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 7748 21428 7800 21480
rect 5448 21360 5500 21412
rect 8024 21360 8076 21412
rect 6736 21292 6788 21344
rect 8760 21292 8812 21344
rect 10784 21632 10836 21684
rect 11888 21632 11940 21684
rect 14004 21632 14056 21684
rect 20260 21632 20312 21684
rect 8944 21428 8996 21480
rect 10508 21496 10560 21548
rect 18052 21564 18104 21616
rect 18144 21564 18196 21616
rect 19248 21564 19300 21616
rect 20904 21564 20956 21616
rect 24400 21564 24452 21616
rect 11612 21496 11664 21548
rect 12808 21496 12860 21548
rect 13636 21496 13688 21548
rect 13176 21428 13228 21480
rect 14096 21496 14148 21548
rect 15568 21496 15620 21548
rect 15844 21496 15896 21548
rect 19340 21539 19392 21548
rect 19340 21505 19349 21539
rect 19349 21505 19383 21539
rect 19383 21505 19392 21539
rect 19340 21496 19392 21505
rect 15108 21428 15160 21480
rect 16396 21428 16448 21480
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 18604 21428 18656 21480
rect 19064 21428 19116 21480
rect 19984 21496 20036 21548
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 22744 21496 22796 21548
rect 23112 21496 23164 21548
rect 24768 21564 24820 21616
rect 30472 21632 30524 21684
rect 30840 21632 30892 21684
rect 31300 21632 31352 21684
rect 26884 21564 26936 21616
rect 26976 21607 27028 21616
rect 26976 21573 26985 21607
rect 26985 21573 27019 21607
rect 27019 21573 27028 21607
rect 26976 21564 27028 21573
rect 27896 21564 27948 21616
rect 21180 21428 21232 21480
rect 22652 21428 22704 21480
rect 25780 21428 25832 21480
rect 25872 21428 25924 21480
rect 26516 21428 26568 21480
rect 26700 21496 26752 21548
rect 28632 21564 28684 21616
rect 30012 21564 30064 21616
rect 30656 21539 30708 21548
rect 30656 21505 30665 21539
rect 30665 21505 30699 21539
rect 30699 21505 30708 21539
rect 30656 21496 30708 21505
rect 31852 21564 31904 21616
rect 10416 21360 10468 21412
rect 10968 21360 11020 21412
rect 14556 21360 14608 21412
rect 16856 21360 16908 21412
rect 19432 21360 19484 21412
rect 23296 21360 23348 21412
rect 25412 21403 25464 21412
rect 25412 21369 25421 21403
rect 25421 21369 25455 21403
rect 25455 21369 25464 21403
rect 25412 21360 25464 21369
rect 26424 21403 26476 21412
rect 26424 21369 26433 21403
rect 26433 21369 26467 21403
rect 26467 21369 26476 21403
rect 28540 21471 28592 21480
rect 26424 21360 26476 21369
rect 13820 21292 13872 21344
rect 14464 21292 14516 21344
rect 16580 21292 16632 21344
rect 18696 21292 18748 21344
rect 20536 21292 20588 21344
rect 21088 21292 21140 21344
rect 23756 21292 23808 21344
rect 24492 21335 24544 21344
rect 24492 21301 24501 21335
rect 24501 21301 24535 21335
rect 24535 21301 24544 21335
rect 24492 21292 24544 21301
rect 26148 21292 26200 21344
rect 28540 21437 28549 21471
rect 28549 21437 28583 21471
rect 28583 21437 28592 21471
rect 28540 21428 28592 21437
rect 28632 21428 28684 21480
rect 29920 21428 29972 21480
rect 32404 21496 32456 21548
rect 33232 21539 33284 21548
rect 29736 21292 29788 21344
rect 31116 21360 31168 21412
rect 33232 21505 33241 21539
rect 33241 21505 33275 21539
rect 33275 21505 33284 21539
rect 33232 21496 33284 21505
rect 33416 21539 33468 21548
rect 33416 21505 33425 21539
rect 33425 21505 33459 21539
rect 33459 21505 33468 21539
rect 33416 21496 33468 21505
rect 34060 21496 34112 21548
rect 34520 21632 34572 21684
rect 35808 21632 35860 21684
rect 34704 21564 34756 21616
rect 36084 21564 36136 21616
rect 37556 21496 37608 21548
rect 33048 21428 33100 21480
rect 34520 21360 34572 21412
rect 31024 21335 31076 21344
rect 31024 21301 31033 21335
rect 31033 21301 31067 21335
rect 31067 21301 31076 21335
rect 31024 21292 31076 21301
rect 32220 21335 32272 21344
rect 32220 21301 32229 21335
rect 32229 21301 32263 21335
rect 32263 21301 32272 21335
rect 32220 21292 32272 21301
rect 34612 21292 34664 21344
rect 37280 21292 37332 21344
rect 37924 21292 37976 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5448 21088 5500 21140
rect 6552 21088 6604 21140
rect 8392 21088 8444 21140
rect 10508 21131 10560 21140
rect 10508 21097 10517 21131
rect 10517 21097 10551 21131
rect 10551 21097 10560 21131
rect 10508 21088 10560 21097
rect 1400 20884 1452 20936
rect 5908 20995 5960 21004
rect 5908 20961 5917 20995
rect 5917 20961 5951 20995
rect 5951 20961 5960 20995
rect 5908 20952 5960 20961
rect 6644 21020 6696 21072
rect 7840 21020 7892 21072
rect 11152 21088 11204 21140
rect 13820 21088 13872 21140
rect 14832 21088 14884 21140
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6000 20884 6052 20893
rect 6460 20884 6512 20936
rect 6736 20884 6788 20936
rect 6000 20748 6052 20800
rect 6736 20748 6788 20800
rect 8116 20884 8168 20936
rect 10784 20952 10836 21004
rect 11152 20995 11204 21004
rect 11152 20961 11161 20995
rect 11161 20961 11195 20995
rect 11195 20961 11204 20995
rect 11152 20952 11204 20961
rect 8300 20859 8352 20868
rect 8300 20825 8309 20859
rect 8309 20825 8343 20859
rect 8343 20825 8352 20859
rect 8300 20816 8352 20825
rect 10968 20927 11020 20936
rect 10968 20893 11003 20927
rect 11003 20893 11020 20927
rect 10968 20884 11020 20893
rect 11336 20816 11388 20868
rect 14004 20952 14056 21004
rect 16396 20952 16448 21004
rect 18236 20952 18288 21004
rect 20076 21088 20128 21140
rect 21180 21131 21232 21140
rect 21180 21097 21189 21131
rect 21189 21097 21223 21131
rect 21223 21097 21232 21131
rect 21180 21088 21232 21097
rect 26240 21088 26292 21140
rect 26332 21088 26384 21140
rect 19432 21020 19484 21072
rect 14740 20884 14792 20936
rect 16580 20884 16632 20936
rect 19340 20884 19392 20936
rect 23572 20952 23624 21004
rect 23848 20952 23900 21004
rect 24584 20952 24636 21004
rect 25504 20952 25556 21004
rect 27712 21020 27764 21072
rect 27896 21131 27948 21140
rect 27896 21097 27905 21131
rect 27905 21097 27939 21131
rect 27939 21097 27948 21131
rect 27896 21088 27948 21097
rect 28172 21088 28224 21140
rect 28540 21088 28592 21140
rect 30012 21131 30064 21140
rect 30012 21097 30021 21131
rect 30021 21097 30055 21131
rect 30055 21097 30064 21131
rect 30012 21088 30064 21097
rect 33416 21088 33468 21140
rect 33692 21131 33744 21140
rect 33692 21097 33701 21131
rect 33701 21097 33735 21131
rect 33735 21097 33744 21131
rect 33692 21088 33744 21097
rect 33784 21088 33836 21140
rect 26884 20952 26936 21004
rect 19984 20884 20036 20936
rect 12808 20816 12860 20868
rect 12900 20816 12952 20868
rect 13544 20816 13596 20868
rect 14648 20816 14700 20868
rect 14924 20816 14976 20868
rect 12440 20791 12492 20800
rect 12440 20757 12449 20791
rect 12449 20757 12483 20791
rect 12483 20757 12492 20791
rect 12440 20748 12492 20757
rect 14004 20748 14056 20800
rect 15568 20748 15620 20800
rect 20904 20884 20956 20936
rect 23204 20884 23256 20936
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 23940 20884 23992 20936
rect 26148 20927 26200 20936
rect 26148 20893 26157 20927
rect 26157 20893 26191 20927
rect 26191 20893 26200 20927
rect 28908 20952 28960 21004
rect 26148 20884 26200 20893
rect 20444 20816 20496 20868
rect 22652 20859 22704 20868
rect 22652 20825 22661 20859
rect 22661 20825 22695 20859
rect 22695 20825 22704 20859
rect 22652 20816 22704 20825
rect 23572 20816 23624 20868
rect 25780 20816 25832 20868
rect 18144 20748 18196 20800
rect 20260 20748 20312 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 26332 20748 26384 20800
rect 27528 20816 27580 20868
rect 26792 20791 26844 20800
rect 26792 20757 26801 20791
rect 26801 20757 26835 20791
rect 26835 20757 26844 20791
rect 26792 20748 26844 20757
rect 28080 20816 28132 20868
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 28908 20816 28960 20868
rect 29092 20816 29144 20868
rect 31116 21020 31168 21072
rect 32036 20952 32088 21004
rect 33048 20952 33100 21004
rect 35716 21020 35768 21072
rect 36452 20995 36504 21004
rect 36452 20961 36461 20995
rect 36461 20961 36495 20995
rect 36495 20961 36504 20995
rect 36452 20952 36504 20961
rect 38108 20995 38160 21004
rect 38108 20961 38117 20995
rect 38117 20961 38151 20995
rect 38151 20961 38160 20995
rect 38108 20952 38160 20961
rect 30840 20884 30892 20936
rect 33140 20884 33192 20936
rect 31944 20816 31996 20868
rect 33416 20816 33468 20868
rect 35348 20859 35400 20868
rect 35348 20825 35357 20859
rect 35357 20825 35391 20859
rect 35391 20825 35400 20859
rect 35348 20816 35400 20825
rect 37280 20816 37332 20868
rect 34704 20748 34756 20800
rect 35900 20748 35952 20800
rect 36728 20748 36780 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6644 20544 6696 20596
rect 6184 20476 6236 20528
rect 11520 20544 11572 20596
rect 13636 20587 13688 20596
rect 13636 20553 13645 20587
rect 13645 20553 13679 20587
rect 13679 20553 13688 20587
rect 13636 20544 13688 20553
rect 14648 20544 14700 20596
rect 15844 20544 15896 20596
rect 18328 20544 18380 20596
rect 19984 20544 20036 20596
rect 22652 20544 22704 20596
rect 6828 20519 6880 20528
rect 6828 20485 6863 20519
rect 6863 20485 6880 20519
rect 6828 20476 6880 20485
rect 7104 20476 7156 20528
rect 8760 20476 8812 20528
rect 9496 20519 9548 20528
rect 9496 20485 9505 20519
rect 9505 20485 9539 20519
rect 9539 20485 9548 20519
rect 9496 20476 9548 20485
rect 10968 20476 11020 20528
rect 11152 20476 11204 20528
rect 12900 20519 12952 20528
rect 12900 20485 12909 20519
rect 12909 20485 12943 20519
rect 12943 20485 12952 20519
rect 12900 20476 12952 20485
rect 13360 20476 13412 20528
rect 14464 20519 14516 20528
rect 14464 20485 14473 20519
rect 14473 20485 14507 20519
rect 14507 20485 14516 20519
rect 14464 20476 14516 20485
rect 15108 20476 15160 20528
rect 15568 20519 15620 20528
rect 15568 20485 15577 20519
rect 15577 20485 15611 20519
rect 15611 20485 15620 20519
rect 15568 20476 15620 20485
rect 16580 20476 16632 20528
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 4528 20408 4580 20460
rect 6644 20451 6696 20460
rect 6644 20417 6653 20451
rect 6653 20417 6687 20451
rect 6687 20417 6696 20451
rect 7840 20451 7892 20460
rect 6644 20408 6696 20417
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8300 20408 8352 20460
rect 6736 20340 6788 20392
rect 8116 20383 8168 20392
rect 8116 20349 8125 20383
rect 8125 20349 8159 20383
rect 8159 20349 8168 20383
rect 8116 20340 8168 20349
rect 9588 20408 9640 20460
rect 10232 20451 10284 20460
rect 10232 20417 10241 20451
rect 10241 20417 10275 20451
rect 10275 20417 10284 20451
rect 10232 20408 10284 20417
rect 11980 20451 12032 20460
rect 11980 20417 11989 20451
rect 11989 20417 12023 20451
rect 12023 20417 12032 20451
rect 11980 20408 12032 20417
rect 10968 20340 11020 20392
rect 11244 20340 11296 20392
rect 12440 20340 12492 20392
rect 10784 20272 10836 20324
rect 14004 20408 14056 20460
rect 15200 20408 15252 20460
rect 18052 20476 18104 20528
rect 19432 20476 19484 20528
rect 14832 20340 14884 20392
rect 17868 20340 17920 20392
rect 19156 20408 19208 20460
rect 19984 20383 20036 20392
rect 19984 20349 19993 20383
rect 19993 20349 20027 20383
rect 20027 20349 20036 20383
rect 19984 20340 20036 20349
rect 20076 20383 20128 20392
rect 20076 20349 20085 20383
rect 20085 20349 20119 20383
rect 20119 20349 20128 20383
rect 20076 20340 20128 20349
rect 20260 20383 20312 20392
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 21824 20408 21876 20460
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 23664 20476 23716 20528
rect 26792 20544 26844 20596
rect 27804 20587 27856 20596
rect 27804 20553 27813 20587
rect 27813 20553 27847 20587
rect 27847 20553 27856 20587
rect 27804 20544 27856 20553
rect 28172 20544 28224 20596
rect 33416 20587 33468 20596
rect 33416 20553 33425 20587
rect 33425 20553 33459 20587
rect 33459 20553 33468 20587
rect 33416 20544 33468 20553
rect 28264 20476 28316 20528
rect 29000 20476 29052 20528
rect 30012 20476 30064 20528
rect 22652 20408 22704 20460
rect 23296 20408 23348 20460
rect 23388 20383 23440 20392
rect 20260 20340 20312 20349
rect 14924 20272 14976 20324
rect 15108 20272 15160 20324
rect 23388 20349 23397 20383
rect 23397 20349 23431 20383
rect 23431 20349 23440 20383
rect 23388 20340 23440 20349
rect 23756 20340 23808 20392
rect 22744 20272 22796 20324
rect 25136 20315 25188 20324
rect 25136 20281 25145 20315
rect 25145 20281 25179 20315
rect 25179 20281 25188 20315
rect 25136 20272 25188 20281
rect 1584 20204 1636 20256
rect 7472 20247 7524 20256
rect 7472 20213 7481 20247
rect 7481 20213 7515 20247
rect 7515 20213 7524 20247
rect 7472 20204 7524 20213
rect 9772 20204 9824 20256
rect 15384 20247 15436 20256
rect 15384 20213 15393 20247
rect 15393 20213 15427 20247
rect 15427 20213 15436 20247
rect 15384 20204 15436 20213
rect 16764 20204 16816 20256
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 18236 20204 18288 20256
rect 19984 20204 20036 20256
rect 20812 20204 20864 20256
rect 23848 20204 23900 20256
rect 25688 20204 25740 20256
rect 26516 20340 26568 20392
rect 27436 20408 27488 20460
rect 27896 20408 27948 20460
rect 28908 20451 28960 20460
rect 28908 20417 28917 20451
rect 28917 20417 28951 20451
rect 28951 20417 28960 20451
rect 28908 20408 28960 20417
rect 27712 20383 27764 20392
rect 27712 20349 27721 20383
rect 27721 20349 27755 20383
rect 27755 20349 27764 20383
rect 27712 20340 27764 20349
rect 27804 20340 27856 20392
rect 28356 20340 28408 20392
rect 26976 20272 27028 20324
rect 29000 20340 29052 20392
rect 32588 20476 32640 20528
rect 33968 20476 34020 20528
rect 30840 20451 30892 20460
rect 30840 20417 30849 20451
rect 30849 20417 30883 20451
rect 30883 20417 30892 20451
rect 30840 20408 30892 20417
rect 31484 20451 31536 20460
rect 31484 20417 31493 20451
rect 31493 20417 31527 20451
rect 31527 20417 31536 20451
rect 31484 20408 31536 20417
rect 31668 20408 31720 20460
rect 33876 20408 33928 20460
rect 34336 20451 34388 20460
rect 34336 20417 34345 20451
rect 34345 20417 34379 20451
rect 34379 20417 34388 20451
rect 34336 20408 34388 20417
rect 34612 20476 34664 20528
rect 36544 20476 36596 20528
rect 37280 20519 37332 20528
rect 37280 20485 37289 20519
rect 37289 20485 37323 20519
rect 37323 20485 37332 20519
rect 37280 20476 37332 20485
rect 37464 20451 37516 20460
rect 37464 20417 37473 20451
rect 37473 20417 37507 20451
rect 37507 20417 37516 20451
rect 37464 20408 37516 20417
rect 27436 20247 27488 20256
rect 27436 20213 27445 20247
rect 27445 20213 27479 20247
rect 27479 20213 27488 20247
rect 27436 20204 27488 20213
rect 29184 20272 29236 20324
rect 29736 20272 29788 20324
rect 30932 20340 30984 20392
rect 32128 20383 32180 20392
rect 32128 20349 32137 20383
rect 32137 20349 32171 20383
rect 32171 20349 32180 20383
rect 32128 20340 32180 20349
rect 31300 20315 31352 20324
rect 31300 20281 31309 20315
rect 31309 20281 31343 20315
rect 31343 20281 31352 20315
rect 31300 20272 31352 20281
rect 31392 20272 31444 20324
rect 35716 20340 35768 20392
rect 28816 20204 28868 20256
rect 30656 20204 30708 20256
rect 30840 20204 30892 20256
rect 34428 20247 34480 20256
rect 34428 20213 34437 20247
rect 34437 20213 34471 20247
rect 34471 20213 34480 20247
rect 34428 20204 34480 20213
rect 34520 20204 34572 20256
rect 35348 20272 35400 20324
rect 37372 20272 37424 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6644 20000 6696 20052
rect 11980 20000 12032 20052
rect 13360 20000 13412 20052
rect 14648 20000 14700 20052
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 15568 20000 15620 20052
rect 16028 20043 16080 20052
rect 16028 20009 16037 20043
rect 16037 20009 16071 20043
rect 16071 20009 16080 20043
rect 16028 20000 16080 20009
rect 16120 20000 16172 20052
rect 16304 20000 16356 20052
rect 18328 20000 18380 20052
rect 18512 20043 18564 20052
rect 18512 20009 18521 20043
rect 18521 20009 18555 20043
rect 18555 20009 18564 20043
rect 18512 20000 18564 20009
rect 20352 20000 20404 20052
rect 23112 20043 23164 20052
rect 23112 20009 23121 20043
rect 23121 20009 23155 20043
rect 23155 20009 23164 20043
rect 23112 20000 23164 20009
rect 27068 20000 27120 20052
rect 27528 20000 27580 20052
rect 28908 20000 28960 20052
rect 30104 20000 30156 20052
rect 31392 20000 31444 20052
rect 32312 20000 32364 20052
rect 35716 20043 35768 20052
rect 35716 20009 35725 20043
rect 35725 20009 35759 20043
rect 35759 20009 35768 20043
rect 35716 20000 35768 20009
rect 6460 19932 6512 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 1584 19907 1636 19916
rect 1584 19873 1593 19907
rect 1593 19873 1627 19907
rect 1627 19873 1636 19907
rect 1584 19864 1636 19873
rect 1860 19907 1912 19916
rect 1860 19873 1869 19907
rect 1869 19873 1903 19907
rect 1903 19873 1912 19907
rect 1860 19864 1912 19873
rect 7104 19907 7156 19916
rect 7104 19873 7113 19907
rect 7113 19873 7147 19907
rect 7147 19873 7156 19907
rect 7104 19864 7156 19873
rect 8116 19864 8168 19916
rect 6736 19796 6788 19848
rect 8668 19796 8720 19848
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 9588 19796 9640 19848
rect 13084 19864 13136 19916
rect 15384 19932 15436 19984
rect 11060 19796 11112 19848
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 13728 19864 13780 19916
rect 14096 19864 14148 19916
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 16672 19932 16724 19984
rect 17316 19932 17368 19984
rect 14556 19864 14608 19873
rect 16764 19864 16816 19916
rect 18236 19864 18288 19916
rect 19340 19932 19392 19984
rect 23204 19932 23256 19984
rect 20720 19907 20772 19916
rect 9036 19728 9088 19780
rect 13084 19728 13136 19780
rect 13544 19728 13596 19780
rect 14648 19796 14700 19848
rect 15200 19728 15252 19780
rect 15844 19796 15896 19848
rect 16580 19796 16632 19848
rect 16856 19839 16908 19848
rect 16856 19805 16865 19839
rect 16865 19805 16899 19839
rect 16899 19805 16908 19839
rect 16856 19796 16908 19805
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 17500 19839 17552 19848
rect 17500 19805 17509 19839
rect 17509 19805 17543 19839
rect 17543 19805 17552 19839
rect 17500 19796 17552 19805
rect 17132 19728 17184 19780
rect 19156 19728 19208 19780
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 10784 19703 10836 19712
rect 10784 19669 10793 19703
rect 10793 19669 10827 19703
rect 10827 19669 10836 19703
rect 10784 19660 10836 19669
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 13452 19703 13504 19712
rect 13452 19669 13461 19703
rect 13461 19669 13495 19703
rect 13495 19669 13504 19703
rect 13452 19660 13504 19669
rect 13820 19660 13872 19712
rect 15108 19660 15160 19712
rect 18328 19660 18380 19712
rect 20720 19873 20729 19907
rect 20729 19873 20763 19907
rect 20763 19873 20772 19907
rect 20720 19864 20772 19873
rect 28356 19864 28408 19916
rect 32496 19932 32548 19984
rect 37832 19932 37884 19984
rect 22376 19839 22428 19848
rect 22376 19805 22385 19839
rect 22385 19805 22419 19839
rect 22419 19805 22428 19839
rect 22376 19796 22428 19805
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 24492 19796 24544 19848
rect 24952 19796 25004 19848
rect 25136 19796 25188 19848
rect 26516 19796 26568 19848
rect 28448 19796 28500 19848
rect 28908 19864 28960 19916
rect 29644 19864 29696 19916
rect 31116 19907 31168 19916
rect 31116 19873 31125 19907
rect 31125 19873 31159 19907
rect 31159 19873 31168 19907
rect 31116 19864 31168 19873
rect 24124 19728 24176 19780
rect 27436 19771 27488 19780
rect 27436 19737 27463 19771
rect 27463 19737 27488 19771
rect 27436 19728 27488 19737
rect 27620 19771 27672 19780
rect 27620 19737 27629 19771
rect 27629 19737 27663 19771
rect 27663 19737 27672 19771
rect 27620 19728 27672 19737
rect 29552 19839 29604 19848
rect 29552 19805 29561 19839
rect 29561 19805 29595 19839
rect 29595 19805 29604 19839
rect 29552 19796 29604 19805
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 20904 19660 20956 19712
rect 23848 19660 23900 19712
rect 27712 19660 27764 19712
rect 29828 19728 29880 19780
rect 30564 19796 30616 19848
rect 30840 19796 30892 19848
rect 32036 19839 32088 19848
rect 32036 19805 32045 19839
rect 32045 19805 32079 19839
rect 32079 19805 32088 19839
rect 32036 19796 32088 19805
rect 32220 19839 32272 19848
rect 32220 19805 32229 19839
rect 32229 19805 32263 19839
rect 32263 19805 32272 19839
rect 32220 19796 32272 19805
rect 31668 19728 31720 19780
rect 32956 19796 33008 19848
rect 34428 19864 34480 19916
rect 37096 19907 37148 19916
rect 33416 19839 33468 19848
rect 33416 19805 33425 19839
rect 33425 19805 33459 19839
rect 33459 19805 33468 19839
rect 33416 19796 33468 19805
rect 34704 19796 34756 19848
rect 34980 19796 35032 19848
rect 37096 19873 37105 19907
rect 37105 19873 37139 19907
rect 37139 19873 37148 19907
rect 37096 19864 37148 19873
rect 37924 19907 37976 19916
rect 37924 19873 37933 19907
rect 37933 19873 37967 19907
rect 37967 19873 37976 19907
rect 37924 19864 37976 19873
rect 35440 19839 35492 19848
rect 35440 19805 35449 19839
rect 35449 19805 35483 19839
rect 35483 19805 35492 19839
rect 35440 19796 35492 19805
rect 35532 19728 35584 19780
rect 30656 19660 30708 19712
rect 30932 19703 30984 19712
rect 30932 19669 30941 19703
rect 30941 19669 30975 19703
rect 30975 19669 30984 19703
rect 30932 19660 30984 19669
rect 33324 19703 33376 19712
rect 33324 19669 33333 19703
rect 33333 19669 33367 19703
rect 33367 19669 33376 19703
rect 33324 19660 33376 19669
rect 33508 19703 33560 19712
rect 33508 19669 33517 19703
rect 33517 19669 33551 19703
rect 33551 19669 33560 19703
rect 33508 19660 33560 19669
rect 33784 19660 33836 19712
rect 34888 19660 34940 19712
rect 37372 19660 37424 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 7104 19456 7156 19508
rect 4620 19320 4672 19372
rect 8668 19388 8720 19440
rect 6460 19320 6512 19372
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 9864 19456 9916 19465
rect 10784 19456 10836 19508
rect 8944 19388 8996 19440
rect 13728 19456 13780 19508
rect 14556 19456 14608 19508
rect 16764 19456 16816 19508
rect 17040 19456 17092 19508
rect 18328 19456 18380 19508
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 2136 19295 2188 19304
rect 2136 19261 2145 19295
rect 2145 19261 2179 19295
rect 2179 19261 2188 19295
rect 2136 19252 2188 19261
rect 9036 19320 9088 19372
rect 11612 19320 11664 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 10324 19252 10376 19304
rect 15200 19388 15252 19440
rect 16396 19388 16448 19440
rect 14188 19320 14240 19372
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 15108 19363 15160 19372
rect 15108 19329 15117 19363
rect 15117 19329 15151 19363
rect 15151 19329 15160 19363
rect 15108 19320 15160 19329
rect 18236 19388 18288 19440
rect 14648 19252 14700 19304
rect 17224 19320 17276 19372
rect 20076 19456 20128 19508
rect 19984 19431 20036 19440
rect 19984 19397 20018 19431
rect 20018 19397 20036 19431
rect 19984 19388 20036 19397
rect 22468 19388 22520 19440
rect 23020 19388 23072 19440
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 23388 19320 23440 19372
rect 25044 19456 25096 19508
rect 26884 19456 26936 19508
rect 27988 19456 28040 19508
rect 28448 19456 28500 19508
rect 28908 19456 28960 19508
rect 29644 19456 29696 19508
rect 30380 19456 30432 19508
rect 31024 19456 31076 19508
rect 33324 19456 33376 19508
rect 33968 19456 34020 19508
rect 24860 19320 24912 19372
rect 25412 19320 25464 19372
rect 18788 19252 18840 19304
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 19432 19252 19484 19304
rect 23020 19252 23072 19304
rect 23756 19295 23808 19304
rect 23756 19261 23765 19295
rect 23765 19261 23799 19295
rect 23799 19261 23808 19295
rect 23756 19252 23808 19261
rect 26056 19252 26108 19304
rect 26976 19320 27028 19372
rect 28264 19363 28316 19372
rect 10232 19184 10284 19236
rect 11152 19184 11204 19236
rect 7840 19116 7892 19168
rect 11796 19116 11848 19168
rect 12808 19116 12860 19168
rect 13084 19116 13136 19168
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 15752 19159 15804 19168
rect 15752 19125 15761 19159
rect 15761 19125 15795 19159
rect 15795 19125 15804 19159
rect 15752 19116 15804 19125
rect 16028 19184 16080 19236
rect 19248 19184 19300 19236
rect 24768 19184 24820 19236
rect 25688 19184 25740 19236
rect 25872 19184 25924 19236
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 28448 19363 28500 19372
rect 28448 19329 28457 19363
rect 28457 19329 28491 19363
rect 28491 19329 28500 19363
rect 28448 19320 28500 19329
rect 29184 19363 29236 19372
rect 29184 19329 29193 19363
rect 29193 19329 29227 19363
rect 29227 19329 29236 19363
rect 29184 19320 29236 19329
rect 28080 19295 28132 19304
rect 28080 19261 28089 19295
rect 28089 19261 28123 19295
rect 28123 19261 28132 19295
rect 28080 19252 28132 19261
rect 29092 19295 29144 19304
rect 29092 19261 29101 19295
rect 29101 19261 29135 19295
rect 29135 19261 29144 19295
rect 29828 19320 29880 19372
rect 30104 19320 30156 19372
rect 32956 19388 33008 19440
rect 33140 19320 33192 19372
rect 33416 19320 33468 19372
rect 29092 19252 29144 19261
rect 18052 19159 18104 19168
rect 18052 19125 18061 19159
rect 18061 19125 18095 19159
rect 18095 19125 18104 19159
rect 18052 19116 18104 19125
rect 20904 19116 20956 19168
rect 21732 19116 21784 19168
rect 22008 19116 22060 19168
rect 22560 19116 22612 19168
rect 23296 19116 23348 19168
rect 25412 19116 25464 19168
rect 25964 19159 26016 19168
rect 25964 19125 25973 19159
rect 25973 19125 26007 19159
rect 26007 19125 26016 19159
rect 25964 19116 26016 19125
rect 28448 19184 28500 19236
rect 30564 19252 30616 19304
rect 31484 19252 31536 19304
rect 31576 19295 31628 19304
rect 31576 19261 31585 19295
rect 31585 19261 31619 19295
rect 31619 19261 31628 19295
rect 31576 19252 31628 19261
rect 32312 19252 32364 19304
rect 34520 19431 34572 19440
rect 34520 19397 34529 19431
rect 34529 19397 34563 19431
rect 34563 19397 34572 19431
rect 34520 19388 34572 19397
rect 36544 19456 36596 19508
rect 36728 19499 36780 19508
rect 36728 19465 36737 19499
rect 36737 19465 36771 19499
rect 36771 19465 36780 19499
rect 36728 19456 36780 19465
rect 35900 19388 35952 19440
rect 37372 19388 37424 19440
rect 37464 19363 37516 19372
rect 34520 19252 34572 19304
rect 34888 19252 34940 19304
rect 35348 19252 35400 19304
rect 35808 19252 35860 19304
rect 37464 19329 37473 19363
rect 37473 19329 37507 19363
rect 37507 19329 37516 19363
rect 37464 19320 37516 19329
rect 30380 19184 30432 19236
rect 26516 19116 26568 19168
rect 30196 19116 30248 19168
rect 32220 19116 32272 19168
rect 32312 19159 32364 19168
rect 32312 19125 32321 19159
rect 32321 19125 32355 19159
rect 32355 19125 32364 19159
rect 32312 19116 32364 19125
rect 32496 19159 32548 19168
rect 32496 19125 32505 19159
rect 32505 19125 32539 19159
rect 32539 19125 32548 19159
rect 32496 19116 32548 19125
rect 33232 19116 33284 19168
rect 34428 19116 34480 19168
rect 35440 19116 35492 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1676 18912 1728 18964
rect 1860 18912 1912 18964
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 14556 18912 14608 18964
rect 15844 18912 15896 18964
rect 10784 18844 10836 18896
rect 9864 18776 9916 18828
rect 10324 18819 10376 18828
rect 10324 18785 10333 18819
rect 10333 18785 10367 18819
rect 10367 18785 10376 18819
rect 10324 18776 10376 18785
rect 2320 18708 2372 18760
rect 7472 18708 7524 18760
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 9680 18708 9732 18760
rect 11888 18776 11940 18828
rect 13912 18844 13964 18896
rect 15200 18844 15252 18896
rect 20352 18912 20404 18964
rect 17684 18844 17736 18896
rect 18696 18844 18748 18896
rect 18788 18844 18840 18896
rect 21364 18844 21416 18896
rect 17224 18776 17276 18828
rect 17500 18776 17552 18828
rect 18236 18776 18288 18828
rect 18512 18776 18564 18828
rect 21548 18776 21600 18828
rect 23664 18912 23716 18964
rect 24216 18912 24268 18964
rect 26240 18955 26292 18964
rect 23388 18844 23440 18896
rect 25872 18844 25924 18896
rect 26240 18921 26249 18955
rect 26249 18921 26283 18955
rect 26283 18921 26292 18955
rect 26240 18912 26292 18921
rect 27988 18955 28040 18964
rect 27988 18921 27997 18955
rect 27997 18921 28031 18955
rect 28031 18921 28040 18955
rect 27988 18912 28040 18921
rect 28540 18844 28592 18896
rect 29276 18912 29328 18964
rect 30104 18844 30156 18896
rect 26332 18819 26384 18828
rect 10692 18708 10744 18760
rect 11796 18708 11848 18760
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 12256 18751 12308 18760
rect 12256 18717 12265 18751
rect 12265 18717 12299 18751
rect 12299 18717 12308 18751
rect 13084 18751 13136 18760
rect 12256 18708 12308 18717
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 15568 18708 15620 18760
rect 16396 18640 16448 18692
rect 17040 18708 17092 18760
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 17316 18640 17368 18692
rect 8300 18572 8352 18624
rect 10508 18572 10560 18624
rect 10784 18572 10836 18624
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 13176 18572 13228 18624
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 15384 18615 15436 18624
rect 13268 18572 13320 18581
rect 15384 18581 15393 18615
rect 15393 18581 15427 18615
rect 15427 18581 15436 18615
rect 15384 18572 15436 18581
rect 16488 18572 16540 18624
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 18604 18708 18656 18760
rect 20812 18708 20864 18760
rect 22100 18708 22152 18760
rect 22928 18751 22980 18760
rect 22928 18717 22937 18751
rect 22937 18717 22971 18751
rect 22971 18717 22980 18751
rect 22928 18708 22980 18717
rect 23296 18708 23348 18760
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 26332 18785 26341 18819
rect 26341 18785 26375 18819
rect 26375 18785 26384 18819
rect 26332 18776 26384 18785
rect 30288 18844 30340 18896
rect 18052 18640 18104 18692
rect 21732 18640 21784 18692
rect 26884 18708 26936 18760
rect 16948 18572 17000 18581
rect 18512 18572 18564 18624
rect 19156 18572 19208 18624
rect 26056 18640 26108 18692
rect 26148 18683 26200 18692
rect 26148 18649 26157 18683
rect 26157 18649 26191 18683
rect 26191 18649 26200 18683
rect 26148 18640 26200 18649
rect 22744 18615 22796 18624
rect 22744 18581 22753 18615
rect 22753 18581 22787 18615
rect 22787 18581 22796 18615
rect 22744 18572 22796 18581
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 25228 18615 25280 18624
rect 25228 18581 25237 18615
rect 25237 18581 25271 18615
rect 25271 18581 25280 18615
rect 25228 18572 25280 18581
rect 26976 18640 27028 18692
rect 29092 18708 29144 18760
rect 27620 18572 27672 18624
rect 28264 18640 28316 18692
rect 29552 18640 29604 18692
rect 30012 18751 30064 18760
rect 30012 18717 30021 18751
rect 30021 18717 30055 18751
rect 30055 18717 30064 18751
rect 30196 18751 30248 18760
rect 30012 18708 30064 18717
rect 30196 18717 30205 18751
rect 30205 18717 30239 18751
rect 30239 18717 30248 18751
rect 30196 18708 30248 18717
rect 30748 18912 30800 18964
rect 30840 18912 30892 18964
rect 31392 18912 31444 18964
rect 31576 18912 31628 18964
rect 34336 18912 34388 18964
rect 35900 18912 35952 18964
rect 31208 18844 31260 18896
rect 35532 18844 35584 18896
rect 36544 18844 36596 18896
rect 35900 18776 35952 18828
rect 31116 18708 31168 18760
rect 31024 18640 31076 18692
rect 32220 18708 32272 18760
rect 33048 18708 33100 18760
rect 32496 18640 32548 18692
rect 33232 18683 33284 18692
rect 33232 18649 33241 18683
rect 33241 18649 33275 18683
rect 33275 18649 33284 18683
rect 33232 18640 33284 18649
rect 33324 18640 33376 18692
rect 29000 18572 29052 18624
rect 30012 18572 30064 18624
rect 31116 18615 31168 18624
rect 31116 18581 31125 18615
rect 31125 18581 31159 18615
rect 31159 18581 31168 18615
rect 31116 18572 31168 18581
rect 32404 18615 32456 18624
rect 32404 18581 32413 18615
rect 32413 18581 32447 18615
rect 32447 18581 32456 18615
rect 32404 18572 32456 18581
rect 33140 18572 33192 18624
rect 33692 18572 33744 18624
rect 34796 18708 34848 18760
rect 35624 18708 35676 18760
rect 35992 18708 36044 18760
rect 34428 18640 34480 18692
rect 34796 18572 34848 18624
rect 34888 18615 34940 18624
rect 34888 18581 34913 18615
rect 34913 18581 34940 18615
rect 34888 18572 34940 18581
rect 35440 18572 35492 18624
rect 36360 18640 36412 18692
rect 37648 18683 37700 18692
rect 37648 18649 37657 18683
rect 37657 18649 37691 18683
rect 37691 18649 37700 18683
rect 37648 18640 37700 18649
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 9588 18368 9640 18420
rect 10784 18411 10836 18420
rect 10784 18377 10793 18411
rect 10793 18377 10827 18411
rect 10827 18377 10836 18411
rect 10784 18368 10836 18377
rect 11612 18368 11664 18420
rect 16948 18368 17000 18420
rect 20076 18368 20128 18420
rect 21548 18368 21600 18420
rect 24952 18411 25004 18420
rect 24952 18377 24961 18411
rect 24961 18377 24995 18411
rect 24995 18377 25004 18411
rect 24952 18368 25004 18377
rect 25964 18411 26016 18420
rect 25964 18377 25991 18411
rect 25991 18377 26016 18411
rect 25964 18368 26016 18377
rect 8668 18300 8720 18352
rect 13268 18300 13320 18352
rect 13452 18300 13504 18352
rect 8300 18275 8352 18284
rect 8300 18241 8334 18275
rect 8334 18241 8352 18275
rect 8300 18232 8352 18241
rect 11612 18232 11664 18284
rect 13820 18232 13872 18284
rect 19340 18300 19392 18352
rect 15752 18232 15804 18284
rect 19248 18275 19300 18284
rect 19248 18241 19266 18275
rect 19266 18241 19300 18275
rect 19248 18232 19300 18241
rect 19432 18232 19484 18284
rect 21364 18300 21416 18352
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 22100 18300 22152 18352
rect 22560 18300 22612 18352
rect 20352 18232 20404 18241
rect 10508 18207 10560 18216
rect 10508 18173 10517 18207
rect 10517 18173 10551 18207
rect 10551 18173 10560 18207
rect 10508 18164 10560 18173
rect 11244 18164 11296 18216
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 12256 18164 12308 18216
rect 13268 18207 13320 18216
rect 12164 18096 12216 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 11428 18028 11480 18080
rect 13268 18173 13277 18207
rect 13277 18173 13311 18207
rect 13311 18173 13320 18207
rect 13268 18164 13320 18173
rect 13912 18164 13964 18216
rect 14924 18164 14976 18216
rect 16580 18164 16632 18216
rect 17040 18164 17092 18216
rect 12808 18096 12860 18148
rect 17224 18139 17276 18148
rect 17224 18105 17233 18139
rect 17233 18105 17267 18139
rect 17267 18105 17276 18139
rect 17224 18096 17276 18105
rect 16580 18028 16632 18080
rect 16764 18028 16816 18080
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 18236 18028 18288 18080
rect 20352 18028 20404 18080
rect 23848 18300 23900 18352
rect 24216 18232 24268 18284
rect 24584 18300 24636 18352
rect 26424 18368 26476 18420
rect 27068 18368 27120 18420
rect 31024 18368 31076 18420
rect 31668 18368 31720 18420
rect 32956 18368 33008 18420
rect 33508 18368 33560 18420
rect 34796 18368 34848 18420
rect 36728 18368 36780 18420
rect 37648 18368 37700 18420
rect 26148 18343 26200 18352
rect 26148 18309 26157 18343
rect 26157 18309 26191 18343
rect 26191 18309 26200 18343
rect 26148 18300 26200 18309
rect 26884 18300 26936 18352
rect 27252 18275 27304 18284
rect 27252 18241 27261 18275
rect 27261 18241 27295 18275
rect 27295 18241 27304 18275
rect 27252 18232 27304 18241
rect 28264 18275 28316 18284
rect 28264 18241 28273 18275
rect 28273 18241 28307 18275
rect 28307 18241 28316 18275
rect 28264 18232 28316 18241
rect 30656 18300 30708 18352
rect 35900 18300 35952 18352
rect 31484 18232 31536 18284
rect 32864 18275 32916 18284
rect 32864 18241 32873 18275
rect 32873 18241 32907 18275
rect 32907 18241 32916 18275
rect 32864 18232 32916 18241
rect 33048 18232 33100 18284
rect 36084 18232 36136 18284
rect 36176 18232 36228 18284
rect 26332 18164 26384 18216
rect 25136 18096 25188 18148
rect 25228 18096 25280 18148
rect 27712 18164 27764 18216
rect 30104 18207 30156 18216
rect 30104 18173 30113 18207
rect 30113 18173 30147 18207
rect 30147 18173 30156 18207
rect 30104 18164 30156 18173
rect 31668 18164 31720 18216
rect 34520 18207 34572 18216
rect 34520 18173 34529 18207
rect 34529 18173 34563 18207
rect 34563 18173 34572 18207
rect 34520 18164 34572 18173
rect 34612 18164 34664 18216
rect 23848 18028 23900 18080
rect 24952 18028 25004 18080
rect 32404 18096 32456 18148
rect 32680 18139 32732 18148
rect 32680 18105 32689 18139
rect 32689 18105 32723 18139
rect 32723 18105 32732 18139
rect 32680 18096 32732 18105
rect 26056 18028 26108 18080
rect 28080 18028 28132 18080
rect 28448 18028 28500 18080
rect 31116 18028 31168 18080
rect 32956 18028 33008 18080
rect 36268 18028 36320 18080
rect 36636 18071 36688 18080
rect 36636 18037 36645 18071
rect 36645 18037 36679 18071
rect 36679 18037 36688 18071
rect 36636 18028 36688 18037
rect 37924 18028 37976 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1676 17688 1728 17740
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 11244 17824 11296 17876
rect 15844 17824 15896 17876
rect 18604 17867 18656 17876
rect 18604 17833 18613 17867
rect 18613 17833 18647 17867
rect 18647 17833 18656 17867
rect 18604 17824 18656 17833
rect 19248 17867 19300 17876
rect 19248 17833 19257 17867
rect 19257 17833 19291 17867
rect 19291 17833 19300 17867
rect 19248 17824 19300 17833
rect 19340 17824 19392 17876
rect 23480 17824 23532 17876
rect 23756 17824 23808 17876
rect 26056 17824 26108 17876
rect 26332 17867 26384 17876
rect 26332 17833 26341 17867
rect 26341 17833 26375 17867
rect 26375 17833 26384 17867
rect 26332 17824 26384 17833
rect 29920 17824 29972 17876
rect 24860 17756 24912 17808
rect 25136 17756 25188 17808
rect 26240 17756 26292 17808
rect 9680 17688 9732 17740
rect 10232 17688 10284 17740
rect 14740 17731 14792 17740
rect 14740 17697 14749 17731
rect 14749 17697 14783 17731
rect 14783 17697 14792 17731
rect 14740 17688 14792 17697
rect 16672 17688 16724 17740
rect 18420 17731 18472 17740
rect 18420 17697 18429 17731
rect 18429 17697 18463 17731
rect 18463 17697 18472 17731
rect 18420 17688 18472 17697
rect 20352 17688 20404 17740
rect 1952 17552 2004 17604
rect 8024 17484 8076 17536
rect 9956 17552 10008 17604
rect 9772 17484 9824 17536
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 11244 17663 11296 17672
rect 10692 17620 10744 17629
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 12164 17620 12216 17672
rect 12992 17620 13044 17672
rect 13360 17620 13412 17672
rect 11612 17552 11664 17604
rect 13912 17552 13964 17604
rect 11520 17484 11572 17536
rect 11796 17484 11848 17536
rect 14556 17620 14608 17672
rect 16580 17620 16632 17672
rect 17224 17620 17276 17672
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 18972 17620 19024 17672
rect 22376 17688 22428 17740
rect 22652 17620 22704 17672
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 23296 17620 23348 17672
rect 23848 17663 23900 17672
rect 23848 17629 23857 17663
rect 23857 17629 23891 17663
rect 23891 17629 23900 17663
rect 23848 17620 23900 17629
rect 24952 17620 25004 17672
rect 15200 17552 15252 17604
rect 16488 17552 16540 17604
rect 23572 17552 23624 17604
rect 15844 17484 15896 17536
rect 20720 17484 20772 17536
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 23848 17484 23900 17536
rect 24584 17484 24636 17536
rect 27620 17688 27672 17740
rect 26884 17620 26936 17672
rect 27528 17620 27580 17672
rect 30656 17756 30708 17808
rect 32864 17824 32916 17876
rect 33048 17824 33100 17876
rect 34520 17824 34572 17876
rect 35348 17824 35400 17876
rect 28724 17688 28776 17740
rect 32772 17756 32824 17808
rect 33876 17756 33928 17808
rect 35256 17756 35308 17808
rect 35440 17756 35492 17808
rect 37464 17756 37516 17808
rect 38016 17756 38068 17808
rect 37096 17731 37148 17740
rect 29828 17620 29880 17672
rect 30104 17620 30156 17672
rect 26516 17484 26568 17536
rect 26700 17527 26752 17536
rect 26700 17493 26709 17527
rect 26709 17493 26743 17527
rect 26743 17493 26752 17527
rect 26700 17484 26752 17493
rect 27712 17552 27764 17604
rect 28264 17552 28316 17604
rect 33232 17620 33284 17672
rect 37096 17697 37105 17731
rect 37105 17697 37139 17731
rect 37139 17697 37148 17731
rect 37096 17688 37148 17697
rect 37924 17731 37976 17740
rect 37924 17697 37933 17731
rect 37933 17697 37967 17731
rect 37967 17697 37976 17731
rect 37924 17688 37976 17697
rect 33692 17620 33744 17672
rect 35256 17620 35308 17672
rect 35532 17620 35584 17672
rect 35808 17620 35860 17672
rect 27160 17484 27212 17536
rect 30748 17484 30800 17536
rect 31392 17484 31444 17536
rect 32956 17552 33008 17604
rect 32404 17484 32456 17536
rect 32496 17527 32548 17536
rect 32496 17493 32521 17527
rect 32521 17493 32548 17527
rect 34888 17527 34940 17536
rect 32496 17484 32548 17493
rect 34888 17493 34897 17527
rect 34897 17493 34931 17527
rect 34931 17493 34940 17527
rect 34888 17484 34940 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 9680 17280 9732 17332
rect 10508 17280 10560 17332
rect 10784 17323 10836 17332
rect 10784 17289 10793 17323
rect 10793 17289 10827 17323
rect 10827 17289 10836 17323
rect 14556 17323 14608 17332
rect 10784 17280 10836 17289
rect 14556 17289 14565 17323
rect 14565 17289 14599 17323
rect 14599 17289 14608 17323
rect 14556 17280 14608 17289
rect 15200 17323 15252 17332
rect 15200 17289 15209 17323
rect 15209 17289 15243 17323
rect 15243 17289 15252 17323
rect 15200 17280 15252 17289
rect 16672 17323 16724 17332
rect 16672 17289 16681 17323
rect 16681 17289 16715 17323
rect 16715 17289 16724 17323
rect 16672 17280 16724 17289
rect 18972 17280 19024 17332
rect 22560 17280 22612 17332
rect 24676 17280 24728 17332
rect 27160 17280 27212 17332
rect 27528 17323 27580 17332
rect 27528 17289 27537 17323
rect 27537 17289 27571 17323
rect 27571 17289 27580 17323
rect 27528 17280 27580 17289
rect 27620 17280 27672 17332
rect 32036 17280 32088 17332
rect 32864 17323 32916 17332
rect 32864 17289 32891 17323
rect 32891 17289 32916 17323
rect 32864 17280 32916 17289
rect 33140 17280 33192 17332
rect 34612 17280 34664 17332
rect 34888 17280 34940 17332
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 8668 17212 8720 17264
rect 14004 17212 14056 17264
rect 8024 17187 8076 17196
rect 8024 17153 8058 17187
rect 8058 17153 8076 17187
rect 8024 17144 8076 17153
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 11244 17144 11296 17196
rect 11612 17144 11664 17196
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 13084 17144 13136 17196
rect 15292 17212 15344 17264
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 18144 17212 18196 17264
rect 18420 17212 18472 17264
rect 16304 17144 16356 17196
rect 16948 17144 17000 17196
rect 17960 17144 18012 17196
rect 18512 17187 18564 17196
rect 9956 17119 10008 17128
rect 9956 17085 9965 17119
rect 9965 17085 9999 17119
rect 9999 17085 10008 17119
rect 9956 17076 10008 17085
rect 10968 17008 11020 17060
rect 13452 17076 13504 17128
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 21180 17212 21232 17264
rect 23848 17212 23900 17264
rect 27252 17212 27304 17264
rect 27436 17212 27488 17264
rect 32680 17212 32732 17264
rect 33048 17255 33100 17264
rect 33048 17221 33057 17255
rect 33057 17221 33091 17255
rect 33091 17221 33100 17255
rect 33048 17212 33100 17221
rect 33600 17212 33652 17264
rect 22376 17187 22428 17196
rect 22376 17153 22385 17187
rect 22385 17153 22419 17187
rect 22419 17153 22428 17187
rect 22376 17144 22428 17153
rect 25044 17144 25096 17196
rect 25504 17187 25556 17196
rect 25504 17153 25513 17187
rect 25513 17153 25547 17187
rect 25547 17153 25556 17187
rect 25504 17144 25556 17153
rect 12900 17008 12952 17060
rect 19432 17076 19484 17128
rect 20168 17076 20220 17128
rect 25688 17187 25740 17196
rect 25688 17153 25697 17187
rect 25697 17153 25731 17187
rect 25731 17153 25740 17187
rect 25688 17144 25740 17153
rect 25872 17187 25924 17196
rect 25872 17153 25881 17187
rect 25881 17153 25915 17187
rect 25915 17153 25924 17187
rect 25872 17144 25924 17153
rect 28264 17187 28316 17196
rect 28264 17153 28273 17187
rect 28273 17153 28307 17187
rect 28307 17153 28316 17187
rect 28264 17144 28316 17153
rect 36268 17144 36320 17196
rect 14832 17008 14884 17060
rect 9404 16940 9456 16992
rect 12624 16940 12676 16992
rect 13728 16983 13780 16992
rect 13728 16949 13737 16983
rect 13737 16949 13771 16983
rect 13771 16949 13780 16983
rect 13728 16940 13780 16949
rect 20904 16940 20956 16992
rect 24584 16940 24636 16992
rect 25872 17008 25924 17060
rect 27620 17076 27672 17128
rect 31116 17119 31168 17128
rect 31116 17085 31125 17119
rect 31125 17085 31159 17119
rect 31159 17085 31168 17119
rect 31116 17076 31168 17085
rect 31668 17076 31720 17128
rect 35716 17076 35768 17128
rect 36728 17119 36780 17128
rect 36728 17085 36737 17119
rect 36737 17085 36771 17119
rect 36771 17085 36780 17119
rect 36728 17076 36780 17085
rect 29644 17051 29696 17060
rect 26700 16940 26752 16992
rect 29644 17017 29653 17051
rect 29653 17017 29687 17051
rect 29687 17017 29696 17051
rect 29644 17008 29696 17017
rect 32404 17008 32456 17060
rect 30748 16940 30800 16992
rect 32128 16940 32180 16992
rect 32956 16940 33008 16992
rect 33692 16983 33744 16992
rect 33692 16949 33701 16983
rect 33701 16949 33735 16983
rect 33735 16949 33744 16983
rect 33692 16940 33744 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 10692 16736 10744 16788
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 19340 16736 19392 16788
rect 22744 16736 22796 16788
rect 25688 16736 25740 16788
rect 27804 16736 27856 16788
rect 8668 16600 8720 16652
rect 11980 16668 12032 16720
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 13084 16668 13136 16720
rect 15752 16668 15804 16720
rect 22376 16711 22428 16720
rect 11704 16600 11756 16609
rect 13268 16600 13320 16652
rect 12624 16532 12676 16584
rect 15844 16575 15896 16584
rect 9220 16507 9272 16516
rect 9220 16473 9254 16507
rect 9254 16473 9272 16507
rect 9220 16464 9272 16473
rect 11980 16464 12032 16516
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 17040 16600 17092 16652
rect 22376 16677 22385 16711
rect 22385 16677 22419 16711
rect 22419 16677 22428 16711
rect 22376 16668 22428 16677
rect 23204 16668 23256 16720
rect 27528 16668 27580 16720
rect 27712 16711 27764 16720
rect 27712 16677 27721 16711
rect 27721 16677 27755 16711
rect 27755 16677 27764 16711
rect 27712 16668 27764 16677
rect 27896 16668 27948 16720
rect 16488 16575 16540 16584
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 16580 16575 16632 16584
rect 16580 16541 16589 16575
rect 16589 16541 16623 16575
rect 16623 16541 16632 16575
rect 16764 16575 16816 16584
rect 16580 16532 16632 16541
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 19432 16600 19484 16652
rect 20260 16643 20312 16652
rect 20260 16609 20269 16643
rect 20269 16609 20303 16643
rect 20303 16609 20312 16643
rect 20260 16600 20312 16609
rect 22100 16600 22152 16652
rect 22468 16600 22520 16652
rect 10784 16396 10836 16448
rect 13176 16396 13228 16448
rect 13912 16396 13964 16448
rect 14188 16396 14240 16448
rect 14464 16507 14516 16516
rect 14464 16473 14473 16507
rect 14473 16473 14507 16507
rect 14507 16473 14516 16507
rect 22192 16532 22244 16584
rect 23204 16575 23256 16584
rect 23204 16541 23213 16575
rect 23213 16541 23247 16575
rect 23247 16541 23256 16575
rect 23204 16532 23256 16541
rect 24584 16575 24636 16584
rect 14464 16464 14516 16473
rect 20536 16464 20588 16516
rect 20720 16464 20772 16516
rect 23112 16464 23164 16516
rect 17960 16396 18012 16448
rect 18144 16439 18196 16448
rect 18144 16405 18153 16439
rect 18153 16405 18187 16439
rect 18187 16405 18196 16439
rect 18144 16396 18196 16405
rect 20076 16396 20128 16448
rect 20444 16396 20496 16448
rect 21088 16396 21140 16448
rect 22928 16396 22980 16448
rect 23296 16396 23348 16448
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 24768 16575 24820 16584
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 25872 16600 25924 16652
rect 26976 16643 27028 16652
rect 26976 16609 26985 16643
rect 26985 16609 27019 16643
rect 27019 16609 27028 16643
rect 28080 16668 28132 16720
rect 29644 16736 29696 16788
rect 30288 16736 30340 16788
rect 32128 16779 32180 16788
rect 32128 16745 32137 16779
rect 32137 16745 32171 16779
rect 32171 16745 32180 16779
rect 32128 16736 32180 16745
rect 33876 16779 33928 16788
rect 33876 16745 33885 16779
rect 33885 16745 33919 16779
rect 33919 16745 33928 16779
rect 33876 16736 33928 16745
rect 34704 16779 34756 16788
rect 34704 16745 34713 16779
rect 34713 16745 34747 16779
rect 34747 16745 34756 16779
rect 34704 16736 34756 16745
rect 35348 16736 35400 16788
rect 29368 16668 29420 16720
rect 26976 16600 27028 16609
rect 25412 16532 25464 16584
rect 26148 16532 26200 16584
rect 28632 16643 28684 16652
rect 28632 16609 28641 16643
rect 28641 16609 28675 16643
rect 28675 16609 28684 16643
rect 28632 16600 28684 16609
rect 29644 16600 29696 16652
rect 27528 16575 27580 16584
rect 27528 16541 27537 16575
rect 27537 16541 27571 16575
rect 27571 16541 27580 16575
rect 27528 16532 27580 16541
rect 24492 16464 24544 16516
rect 27712 16464 27764 16516
rect 29184 16532 29236 16584
rect 30196 16668 30248 16720
rect 31944 16711 31996 16720
rect 31944 16677 31953 16711
rect 31953 16677 31987 16711
rect 31987 16677 31996 16711
rect 31944 16668 31996 16677
rect 37464 16668 37516 16720
rect 29644 16464 29696 16516
rect 30380 16464 30432 16516
rect 30932 16532 30984 16584
rect 31484 16575 31536 16584
rect 31484 16541 31493 16575
rect 31493 16541 31527 16575
rect 31527 16541 31536 16575
rect 31484 16532 31536 16541
rect 32772 16575 32824 16584
rect 31024 16464 31076 16516
rect 32220 16464 32272 16516
rect 32772 16541 32781 16575
rect 32781 16541 32815 16575
rect 32815 16541 32824 16575
rect 32772 16532 32824 16541
rect 33048 16575 33100 16584
rect 33048 16541 33057 16575
rect 33057 16541 33091 16575
rect 33091 16541 33100 16575
rect 34704 16600 34756 16652
rect 35348 16600 35400 16652
rect 33048 16532 33100 16541
rect 34520 16532 34572 16584
rect 35900 16600 35952 16652
rect 33324 16464 33376 16516
rect 33692 16507 33744 16516
rect 33692 16473 33701 16507
rect 33701 16473 33735 16507
rect 33735 16473 33744 16507
rect 33692 16464 33744 16473
rect 36268 16464 36320 16516
rect 37924 16464 37976 16516
rect 38108 16507 38160 16516
rect 38108 16473 38117 16507
rect 38117 16473 38151 16507
rect 38151 16473 38160 16507
rect 38108 16464 38160 16473
rect 24860 16396 24912 16448
rect 25504 16396 25556 16448
rect 25780 16396 25832 16448
rect 28080 16396 28132 16448
rect 28264 16396 28316 16448
rect 29736 16396 29788 16448
rect 30104 16396 30156 16448
rect 30472 16396 30524 16448
rect 30748 16439 30800 16448
rect 30748 16405 30757 16439
rect 30757 16405 30791 16439
rect 30791 16405 30800 16439
rect 30748 16396 30800 16405
rect 32496 16396 32548 16448
rect 34796 16396 34848 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 12900 16235 12952 16244
rect 12900 16201 12909 16235
rect 12909 16201 12943 16235
rect 12943 16201 12952 16235
rect 12900 16192 12952 16201
rect 14188 16192 14240 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 20444 16192 20496 16244
rect 23020 16192 23072 16244
rect 27620 16192 27672 16244
rect 29644 16235 29696 16244
rect 29644 16201 29653 16235
rect 29653 16201 29687 16235
rect 29687 16201 29696 16235
rect 29644 16192 29696 16201
rect 31116 16192 31168 16244
rect 34796 16192 34848 16244
rect 8668 16124 8720 16176
rect 12624 16124 12676 16176
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 10968 16056 11020 16108
rect 14740 16124 14792 16176
rect 18144 16124 18196 16176
rect 20628 16124 20680 16176
rect 13912 16099 13964 16108
rect 13912 16065 13946 16099
rect 13946 16065 13964 16099
rect 3240 15852 3292 15904
rect 13912 16056 13964 16065
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 17132 16099 17184 16108
rect 17132 16065 17141 16099
rect 17141 16065 17175 16099
rect 17175 16065 17184 16099
rect 17132 16056 17184 16065
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 23204 16124 23256 16176
rect 24860 16124 24912 16176
rect 25044 16124 25096 16176
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 23112 16099 23164 16108
rect 23112 16065 23121 16099
rect 23121 16065 23155 16099
rect 23155 16065 23164 16099
rect 23112 16056 23164 16065
rect 24216 16099 24268 16108
rect 24216 16065 24225 16099
rect 24225 16065 24259 16099
rect 24259 16065 24268 16099
rect 24216 16056 24268 16065
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 26700 16056 26752 16108
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27252 16056 27304 16108
rect 27620 16056 27672 16108
rect 28080 16124 28132 16176
rect 33140 16124 33192 16176
rect 33876 16124 33928 16176
rect 34520 16124 34572 16176
rect 35532 16124 35584 16176
rect 37924 16192 37976 16244
rect 30748 16056 30800 16108
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 32956 16056 33008 16108
rect 34060 16099 34112 16108
rect 34060 16065 34069 16099
rect 34069 16065 34103 16099
rect 34103 16065 34112 16099
rect 34060 16056 34112 16065
rect 34796 16056 34848 16108
rect 37464 16099 37516 16108
rect 37464 16065 37473 16099
rect 37473 16065 37507 16099
rect 37507 16065 37516 16099
rect 37464 16056 37516 16065
rect 37832 16056 37884 16108
rect 12716 15852 12768 15904
rect 15844 15895 15896 15904
rect 15844 15861 15853 15895
rect 15853 15861 15887 15895
rect 15887 15861 15896 15895
rect 15844 15852 15896 15861
rect 16672 15852 16724 15904
rect 17868 15988 17920 16040
rect 18236 16031 18288 16040
rect 18236 15997 18245 16031
rect 18245 15997 18279 16031
rect 18279 15997 18288 16031
rect 18236 15988 18288 15997
rect 20536 15920 20588 15972
rect 24492 15988 24544 16040
rect 30288 16031 30340 16040
rect 30288 15997 30297 16031
rect 30297 15997 30331 16031
rect 30331 15997 30340 16031
rect 30288 15988 30340 15997
rect 19800 15852 19852 15904
rect 21548 15852 21600 15904
rect 27436 15920 27488 15972
rect 29184 15920 29236 15972
rect 30472 15920 30524 15972
rect 32588 15988 32640 16040
rect 36544 16031 36596 16040
rect 36544 15997 36553 16031
rect 36553 15997 36587 16031
rect 36587 15997 36596 16031
rect 36544 15988 36596 15997
rect 22928 15895 22980 15904
rect 22928 15861 22937 15895
rect 22937 15861 22971 15895
rect 22971 15861 22980 15895
rect 22928 15852 22980 15861
rect 25504 15852 25556 15904
rect 27988 15852 28040 15904
rect 28356 15852 28408 15904
rect 31668 15852 31720 15904
rect 32956 15895 33008 15904
rect 32956 15861 32965 15895
rect 32965 15861 32999 15895
rect 32999 15861 33008 15895
rect 32956 15852 33008 15861
rect 33324 15852 33376 15904
rect 34336 15895 34388 15904
rect 34336 15861 34345 15895
rect 34345 15861 34379 15895
rect 34379 15861 34388 15895
rect 34336 15852 34388 15861
rect 34704 15920 34756 15972
rect 35716 15852 35768 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 10968 15691 11020 15700
rect 10968 15657 10977 15691
rect 10977 15657 11011 15691
rect 11011 15657 11020 15691
rect 10968 15648 11020 15657
rect 13084 15648 13136 15700
rect 13636 15648 13688 15700
rect 18236 15648 18288 15700
rect 18880 15648 18932 15700
rect 28080 15648 28132 15700
rect 28356 15648 28408 15700
rect 33140 15648 33192 15700
rect 34796 15648 34848 15700
rect 9956 15580 10008 15632
rect 13912 15580 13964 15632
rect 14740 15580 14792 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3240 15555 3292 15564
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 11888 15444 11940 15496
rect 12716 15444 12768 15496
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 20444 15580 20496 15632
rect 22008 15580 22060 15632
rect 22560 15580 22612 15632
rect 23204 15580 23256 15632
rect 26700 15580 26752 15632
rect 19800 15555 19852 15564
rect 19800 15521 19809 15555
rect 19809 15521 19843 15555
rect 19843 15521 19852 15555
rect 19800 15512 19852 15521
rect 21088 15512 21140 15564
rect 25044 15512 25096 15564
rect 25504 15555 25556 15564
rect 25504 15521 25513 15555
rect 25513 15521 25547 15555
rect 25547 15521 25556 15555
rect 25504 15512 25556 15521
rect 27988 15555 28040 15564
rect 27988 15521 27997 15555
rect 27997 15521 28031 15555
rect 28031 15521 28040 15555
rect 27988 15512 28040 15521
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 21824 15444 21876 15496
rect 22192 15444 22244 15496
rect 24952 15444 25004 15496
rect 27804 15444 27856 15496
rect 28264 15487 28316 15496
rect 28264 15453 28273 15487
rect 28273 15453 28307 15487
rect 28307 15453 28316 15487
rect 28264 15444 28316 15453
rect 32312 15580 32364 15632
rect 30196 15555 30248 15564
rect 30196 15521 30205 15555
rect 30205 15521 30239 15555
rect 30239 15521 30248 15555
rect 30196 15512 30248 15521
rect 31668 15512 31720 15564
rect 34336 15512 34388 15564
rect 35256 15555 35308 15564
rect 35256 15521 35265 15555
rect 35265 15521 35299 15555
rect 35299 15521 35308 15555
rect 35256 15512 35308 15521
rect 37096 15555 37148 15564
rect 37096 15521 37105 15555
rect 37105 15521 37139 15555
rect 37139 15521 37148 15555
rect 37096 15512 37148 15521
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 30380 15487 30432 15496
rect 30380 15453 30389 15487
rect 30389 15453 30423 15487
rect 30423 15453 30432 15487
rect 30380 15444 30432 15453
rect 30472 15487 30524 15496
rect 30472 15453 30481 15487
rect 30481 15453 30515 15487
rect 30515 15453 30524 15487
rect 30472 15444 30524 15453
rect 31208 15444 31260 15496
rect 31484 15444 31536 15496
rect 34060 15444 34112 15496
rect 35440 15487 35492 15496
rect 35440 15453 35449 15487
rect 35449 15453 35483 15487
rect 35483 15453 35492 15487
rect 35440 15444 35492 15453
rect 35624 15444 35676 15496
rect 38108 15487 38160 15496
rect 38108 15453 38117 15487
rect 38117 15453 38151 15487
rect 38151 15453 38160 15487
rect 38108 15444 38160 15453
rect 3056 15419 3108 15428
rect 3056 15385 3065 15419
rect 3065 15385 3099 15419
rect 3099 15385 3108 15419
rect 3056 15376 3108 15385
rect 12532 15376 12584 15428
rect 12624 15376 12676 15428
rect 15108 15419 15160 15428
rect 15108 15385 15117 15419
rect 15117 15385 15151 15419
rect 15151 15385 15160 15419
rect 15108 15376 15160 15385
rect 15844 15376 15896 15428
rect 21548 15419 21600 15428
rect 21548 15385 21557 15419
rect 21557 15385 21591 15419
rect 21591 15385 21600 15419
rect 21548 15376 21600 15385
rect 22008 15376 22060 15428
rect 17500 15351 17552 15360
rect 17500 15317 17509 15351
rect 17509 15317 17543 15351
rect 17543 15317 17552 15351
rect 17500 15308 17552 15317
rect 19432 15308 19484 15360
rect 19984 15308 20036 15360
rect 20536 15308 20588 15360
rect 20904 15308 20956 15360
rect 26424 15308 26476 15360
rect 26884 15308 26936 15360
rect 30564 15351 30616 15360
rect 30564 15317 30573 15351
rect 30573 15317 30607 15351
rect 30607 15317 30616 15351
rect 34704 15376 34756 15428
rect 37924 15419 37976 15428
rect 37924 15385 37933 15419
rect 37933 15385 37967 15419
rect 37967 15385 37976 15419
rect 37924 15376 37976 15385
rect 30564 15308 30616 15317
rect 34520 15308 34572 15360
rect 34796 15308 34848 15360
rect 35256 15308 35308 15360
rect 35716 15308 35768 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 3056 15104 3108 15156
rect 14464 15104 14516 15156
rect 15108 15147 15160 15156
rect 15108 15113 15117 15147
rect 15117 15113 15151 15147
rect 15151 15113 15160 15147
rect 15108 15104 15160 15113
rect 17684 15104 17736 15156
rect 20260 15104 20312 15156
rect 20996 15104 21048 15156
rect 22284 15104 22336 15156
rect 12624 15079 12676 15088
rect 12624 15045 12633 15079
rect 12633 15045 12667 15079
rect 12667 15045 12676 15079
rect 12624 15036 12676 15045
rect 14004 15036 14056 15088
rect 17960 15036 18012 15088
rect 18880 15079 18932 15088
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 7656 14968 7708 15020
rect 13820 14968 13872 15020
rect 15200 15011 15252 15020
rect 12716 14900 12768 14952
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 15200 14968 15252 14977
rect 15568 14968 15620 15020
rect 15752 14900 15804 14952
rect 13636 14875 13688 14884
rect 13636 14841 13645 14875
rect 13645 14841 13679 14875
rect 13679 14841 13688 14875
rect 13636 14832 13688 14841
rect 1860 14807 1912 14816
rect 1860 14773 1869 14807
rect 1869 14773 1903 14807
rect 1903 14773 1912 14807
rect 1860 14764 1912 14773
rect 3056 14764 3108 14816
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 14464 14764 14516 14773
rect 16672 14943 16724 14952
rect 16672 14909 16681 14943
rect 16681 14909 16715 14943
rect 16715 14909 16724 14943
rect 16672 14900 16724 14909
rect 17316 14900 17368 14952
rect 17960 14900 18012 14952
rect 18880 15045 18889 15079
rect 18889 15045 18923 15079
rect 18923 15045 18932 15079
rect 18880 15036 18932 15045
rect 20904 15079 20956 15088
rect 20904 15045 20913 15079
rect 20913 15045 20947 15079
rect 20947 15045 20956 15079
rect 20904 15036 20956 15045
rect 19432 14968 19484 15020
rect 19892 15011 19944 15020
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 20076 14900 20128 14952
rect 21916 14968 21968 15020
rect 23572 15104 23624 15156
rect 25044 15104 25096 15156
rect 25872 15104 25924 15156
rect 29368 15147 29420 15156
rect 29368 15113 29377 15147
rect 29377 15113 29411 15147
rect 29411 15113 29420 15147
rect 29368 15104 29420 15113
rect 29828 15147 29880 15156
rect 29828 15113 29837 15147
rect 29837 15113 29871 15147
rect 29871 15113 29880 15147
rect 29828 15104 29880 15113
rect 30288 15104 30340 15156
rect 26976 15036 27028 15088
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 24860 15011 24912 15020
rect 21824 14943 21876 14952
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 19340 14764 19392 14816
rect 19708 14807 19760 14816
rect 19708 14773 19717 14807
rect 19717 14773 19751 14807
rect 19751 14773 19760 14807
rect 19708 14764 19760 14773
rect 19984 14764 20036 14816
rect 21824 14909 21833 14943
rect 21833 14909 21867 14943
rect 21867 14909 21876 14943
rect 21824 14900 21876 14909
rect 22008 14900 22060 14952
rect 24860 14977 24869 15011
rect 24869 14977 24903 15011
rect 24903 14977 24912 15011
rect 24860 14968 24912 14977
rect 21732 14832 21784 14884
rect 25228 14832 25280 14884
rect 25320 14832 25372 14884
rect 25596 14968 25648 15020
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 26424 14968 26476 14977
rect 29000 15036 29052 15088
rect 31484 15104 31536 15156
rect 32404 15104 32456 15156
rect 31024 15079 31076 15088
rect 26700 14900 26752 14952
rect 27896 14968 27948 15020
rect 27804 14900 27856 14952
rect 29092 14968 29144 15020
rect 31024 15045 31046 15079
rect 31046 15045 31076 15079
rect 31024 15036 31076 15045
rect 31208 15079 31260 15088
rect 31208 15045 31217 15079
rect 31217 15045 31251 15079
rect 31251 15045 31260 15079
rect 31208 15036 31260 15045
rect 32496 15079 32548 15088
rect 32496 15045 32505 15079
rect 32505 15045 32539 15079
rect 32539 15045 32548 15079
rect 32496 15036 32548 15045
rect 29552 14968 29604 15020
rect 30840 14968 30892 15020
rect 31116 14968 31168 15020
rect 31668 14968 31720 15020
rect 36544 15104 36596 15156
rect 33324 15079 33376 15088
rect 33324 15045 33333 15079
rect 33333 15045 33367 15079
rect 33367 15045 33376 15079
rect 33324 15036 33376 15045
rect 34796 15036 34848 15088
rect 35624 15036 35676 15088
rect 36360 15036 36412 15088
rect 34428 14968 34480 15020
rect 35440 15011 35492 15020
rect 35440 14977 35449 15011
rect 35449 14977 35483 15011
rect 35483 14977 35492 15011
rect 35440 14968 35492 14977
rect 35716 15011 35768 15020
rect 35716 14977 35725 15011
rect 35725 14977 35759 15011
rect 35759 14977 35768 15011
rect 35716 14968 35768 14977
rect 35808 14968 35860 15020
rect 38292 14968 38344 15020
rect 31484 14900 31536 14952
rect 32220 14900 32272 14952
rect 35348 14900 35400 14952
rect 21364 14764 21416 14816
rect 21548 14764 21600 14816
rect 25872 14764 25924 14816
rect 29000 14764 29052 14816
rect 35256 14832 35308 14884
rect 30564 14764 30616 14816
rect 31024 14807 31076 14816
rect 31024 14773 31033 14807
rect 31033 14773 31067 14807
rect 31067 14773 31076 14807
rect 31024 14764 31076 14773
rect 32312 14807 32364 14816
rect 32312 14773 32321 14807
rect 32321 14773 32355 14807
rect 32355 14773 32364 14807
rect 32312 14764 32364 14773
rect 32404 14764 32456 14816
rect 33784 14764 33836 14816
rect 35348 14764 35400 14816
rect 35808 14764 35860 14816
rect 36728 14764 36780 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 12532 14560 12584 14612
rect 17316 14603 17368 14612
rect 17316 14569 17325 14603
rect 17325 14569 17359 14603
rect 17359 14569 17368 14603
rect 17316 14560 17368 14569
rect 17500 14560 17552 14612
rect 17868 14560 17920 14612
rect 19064 14560 19116 14612
rect 2780 14492 2832 14544
rect 14556 14492 14608 14544
rect 17224 14492 17276 14544
rect 20904 14560 20956 14612
rect 21732 14560 21784 14612
rect 23296 14560 23348 14612
rect 25412 14560 25464 14612
rect 32312 14560 32364 14612
rect 33876 14560 33928 14612
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 19340 14492 19392 14544
rect 20628 14492 20680 14544
rect 20720 14492 20772 14544
rect 21548 14492 21600 14544
rect 24860 14492 24912 14544
rect 30748 14492 30800 14544
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 15660 14356 15712 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 17040 14356 17092 14408
rect 19708 14424 19760 14476
rect 20812 14424 20864 14476
rect 17960 14356 18012 14408
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 17684 14288 17736 14340
rect 18052 14288 18104 14340
rect 18512 14356 18564 14408
rect 18788 14356 18840 14408
rect 18972 14288 19024 14340
rect 14188 14220 14240 14272
rect 16580 14220 16632 14272
rect 17868 14220 17920 14272
rect 17960 14220 18012 14272
rect 19432 14220 19484 14272
rect 21824 14356 21876 14408
rect 22560 14467 22612 14476
rect 22560 14433 22569 14467
rect 22569 14433 22603 14467
rect 22603 14433 22612 14467
rect 22560 14424 22612 14433
rect 20996 14220 21048 14272
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 21732 14288 21784 14340
rect 22100 14331 22152 14340
rect 22100 14297 22109 14331
rect 22109 14297 22143 14331
rect 22143 14297 22152 14331
rect 23296 14424 23348 14476
rect 23572 14467 23624 14476
rect 23572 14433 23581 14467
rect 23581 14433 23615 14467
rect 23615 14433 23624 14467
rect 23572 14424 23624 14433
rect 25136 14424 25188 14476
rect 29552 14467 29604 14476
rect 29552 14433 29561 14467
rect 29561 14433 29595 14467
rect 29595 14433 29604 14467
rect 29552 14424 29604 14433
rect 30288 14424 30340 14476
rect 31484 14424 31536 14476
rect 31760 14492 31812 14544
rect 37464 14560 37516 14612
rect 34612 14492 34664 14544
rect 35348 14535 35400 14544
rect 35348 14501 35357 14535
rect 35357 14501 35391 14535
rect 35391 14501 35400 14535
rect 35348 14492 35400 14501
rect 22100 14288 22152 14297
rect 30840 14356 30892 14408
rect 31208 14356 31260 14408
rect 32036 14356 32088 14408
rect 36728 14424 36780 14476
rect 38108 14467 38160 14476
rect 38108 14433 38117 14467
rect 38117 14433 38151 14467
rect 38151 14433 38160 14467
rect 38108 14424 38160 14433
rect 23664 14288 23716 14340
rect 25872 14331 25924 14340
rect 25872 14297 25881 14331
rect 25881 14297 25915 14331
rect 25915 14297 25924 14331
rect 25872 14288 25924 14297
rect 23388 14220 23440 14272
rect 27436 14288 27488 14340
rect 32220 14288 32272 14340
rect 34152 14356 34204 14408
rect 36176 14356 36228 14408
rect 33968 14331 34020 14340
rect 33968 14297 33977 14331
rect 33977 14297 34011 14331
rect 34011 14297 34020 14331
rect 35164 14331 35216 14340
rect 33968 14288 34020 14297
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 28816 14220 28868 14272
rect 31576 14220 31628 14272
rect 33600 14263 33652 14272
rect 33600 14229 33609 14263
rect 33609 14229 33643 14263
rect 33643 14229 33652 14263
rect 33600 14220 33652 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 14004 14016 14056 14068
rect 15200 14016 15252 14068
rect 14280 13948 14332 14000
rect 14464 13948 14516 14000
rect 17224 13991 17276 14000
rect 17224 13957 17233 13991
rect 17233 13957 17267 13991
rect 17267 13957 17276 13991
rect 17224 13948 17276 13957
rect 17500 13948 17552 14000
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 19340 14016 19392 14068
rect 21916 14016 21968 14068
rect 18420 13923 18472 13932
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 13820 13812 13872 13864
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 14556 13812 14608 13864
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 20812 13948 20864 14000
rect 21824 13991 21876 14000
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 20168 13880 20220 13932
rect 20444 13880 20496 13932
rect 15936 13812 15988 13864
rect 16764 13812 16816 13864
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 19064 13812 19116 13864
rect 20720 13923 20772 13932
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 20720 13880 20772 13889
rect 21824 13957 21833 13991
rect 21833 13957 21867 13991
rect 21867 13957 21876 13991
rect 21824 13948 21876 13957
rect 21732 13880 21784 13932
rect 22008 13880 22060 13932
rect 25044 14016 25096 14068
rect 25320 14059 25372 14068
rect 25320 14025 25329 14059
rect 25329 14025 25363 14059
rect 25363 14025 25372 14059
rect 25320 14016 25372 14025
rect 27896 14016 27948 14068
rect 29552 14016 29604 14068
rect 30564 14016 30616 14068
rect 31024 14059 31076 14068
rect 31024 14025 31033 14059
rect 31033 14025 31067 14059
rect 31067 14025 31076 14059
rect 31024 14016 31076 14025
rect 31208 14016 31260 14068
rect 35716 14016 35768 14068
rect 37924 14016 37976 14068
rect 26700 13948 26752 14000
rect 27344 13948 27396 14000
rect 28632 13948 28684 14000
rect 25504 13923 25556 13932
rect 25504 13889 25513 13923
rect 25513 13889 25547 13923
rect 25547 13889 25556 13923
rect 25504 13880 25556 13889
rect 26148 13923 26200 13932
rect 26148 13889 26157 13923
rect 26157 13889 26191 13923
rect 26191 13889 26200 13923
rect 26148 13880 26200 13889
rect 26240 13880 26292 13932
rect 31116 13948 31168 14000
rect 31208 13923 31260 13932
rect 31208 13889 31217 13923
rect 31217 13889 31251 13923
rect 31251 13889 31260 13923
rect 31208 13880 31260 13889
rect 31576 13948 31628 14000
rect 20812 13812 20864 13864
rect 23204 13855 23256 13864
rect 5080 13744 5132 13796
rect 10416 13744 10468 13796
rect 17316 13744 17368 13796
rect 19340 13744 19392 13796
rect 19984 13744 20036 13796
rect 21824 13744 21876 13796
rect 15476 13676 15528 13728
rect 19248 13676 19300 13728
rect 20444 13719 20496 13728
rect 20444 13685 20453 13719
rect 20453 13685 20487 13719
rect 20487 13685 20496 13719
rect 20444 13676 20496 13685
rect 20628 13719 20680 13728
rect 20628 13685 20637 13719
rect 20637 13685 20671 13719
rect 20671 13685 20680 13719
rect 20628 13676 20680 13685
rect 21364 13676 21416 13728
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 23296 13812 23348 13864
rect 28632 13812 28684 13864
rect 29368 13812 29420 13864
rect 29920 13855 29972 13864
rect 29920 13821 29929 13855
rect 29929 13821 29963 13855
rect 29963 13821 29972 13855
rect 29920 13812 29972 13821
rect 31116 13812 31168 13864
rect 32036 13880 32088 13932
rect 32956 13880 33008 13932
rect 31576 13855 31628 13864
rect 31576 13821 31585 13855
rect 31585 13821 31619 13855
rect 31619 13821 31628 13855
rect 31576 13812 31628 13821
rect 33232 13880 33284 13932
rect 35440 13948 35492 14000
rect 36544 13948 36596 14000
rect 34152 13923 34204 13932
rect 34152 13889 34161 13923
rect 34161 13889 34195 13923
rect 34195 13889 34204 13923
rect 34152 13880 34204 13889
rect 37464 13923 37516 13932
rect 37464 13889 37473 13923
rect 37473 13889 37507 13923
rect 37507 13889 37516 13923
rect 37464 13880 37516 13889
rect 33876 13855 33928 13864
rect 33876 13821 33885 13855
rect 33885 13821 33919 13855
rect 33919 13821 33928 13855
rect 33876 13812 33928 13821
rect 35716 13812 35768 13864
rect 36452 13855 36504 13864
rect 36452 13821 36461 13855
rect 36461 13821 36495 13855
rect 36495 13821 36504 13855
rect 36452 13812 36504 13821
rect 24768 13676 24820 13728
rect 27160 13676 27212 13728
rect 27988 13676 28040 13728
rect 29552 13676 29604 13728
rect 32588 13676 32640 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2044 13472 2096 13524
rect 4068 13472 4120 13524
rect 15476 13472 15528 13524
rect 15660 13472 15712 13524
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 20352 13515 20404 13524
rect 20352 13481 20361 13515
rect 20361 13481 20395 13515
rect 20395 13481 20404 13515
rect 20352 13472 20404 13481
rect 21088 13472 21140 13524
rect 23204 13515 23256 13524
rect 23204 13481 23213 13515
rect 23213 13481 23247 13515
rect 23247 13481 23256 13515
rect 23204 13472 23256 13481
rect 26240 13472 26292 13524
rect 27896 13472 27948 13524
rect 28540 13472 28592 13524
rect 29644 13515 29696 13524
rect 29644 13481 29653 13515
rect 29653 13481 29687 13515
rect 29687 13481 29696 13515
rect 29644 13472 29696 13481
rect 16672 13336 16724 13388
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 17500 13379 17552 13388
rect 17500 13345 17509 13379
rect 17509 13345 17543 13379
rect 17543 13345 17552 13379
rect 17500 13336 17552 13345
rect 1400 13268 1452 13320
rect 5080 13268 5132 13320
rect 16580 13268 16632 13320
rect 20628 13404 20680 13456
rect 25596 13404 25648 13456
rect 26516 13404 26568 13456
rect 26884 13404 26936 13456
rect 20996 13379 21048 13388
rect 20996 13345 21005 13379
rect 21005 13345 21039 13379
rect 21039 13345 21048 13379
rect 20996 13336 21048 13345
rect 21732 13336 21784 13388
rect 21824 13336 21876 13388
rect 20352 13268 20404 13320
rect 22376 13268 22428 13320
rect 22560 13268 22612 13320
rect 23388 13311 23440 13320
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 24952 13268 25004 13320
rect 14004 13200 14056 13252
rect 16120 13243 16172 13252
rect 16120 13209 16129 13243
rect 16129 13209 16163 13243
rect 16163 13209 16172 13243
rect 16120 13200 16172 13209
rect 18236 13243 18288 13252
rect 18236 13209 18245 13243
rect 18245 13209 18279 13243
rect 18279 13209 18288 13243
rect 18236 13200 18288 13209
rect 20996 13200 21048 13252
rect 21548 13243 21600 13252
rect 21548 13209 21557 13243
rect 21557 13209 21591 13243
rect 21591 13209 21600 13243
rect 21548 13200 21600 13209
rect 21916 13200 21968 13252
rect 22100 13200 22152 13252
rect 23020 13200 23072 13252
rect 23296 13200 23348 13252
rect 23480 13200 23532 13252
rect 25504 13200 25556 13252
rect 25780 13268 25832 13320
rect 26884 13311 26936 13320
rect 26884 13277 26893 13311
rect 26893 13277 26927 13311
rect 26927 13277 26936 13311
rect 26884 13268 26936 13277
rect 16764 13132 16816 13184
rect 18328 13175 18380 13184
rect 18328 13141 18337 13175
rect 18337 13141 18371 13175
rect 18371 13141 18380 13175
rect 18328 13132 18380 13141
rect 19984 13132 20036 13184
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 22192 13132 22244 13184
rect 22468 13132 22520 13184
rect 24308 13132 24360 13184
rect 24768 13132 24820 13184
rect 25688 13175 25740 13184
rect 25688 13141 25697 13175
rect 25697 13141 25731 13175
rect 25731 13141 25740 13175
rect 25688 13132 25740 13141
rect 26056 13132 26108 13184
rect 26332 13175 26384 13184
rect 26332 13141 26341 13175
rect 26341 13141 26375 13175
rect 26375 13141 26384 13175
rect 26332 13132 26384 13141
rect 27068 13175 27120 13184
rect 27068 13141 27077 13175
rect 27077 13141 27111 13175
rect 27111 13141 27120 13175
rect 27068 13132 27120 13141
rect 29276 13336 29328 13388
rect 29460 13336 29512 13388
rect 29920 13472 29972 13524
rect 30656 13472 30708 13524
rect 34152 13515 34204 13524
rect 34152 13481 34161 13515
rect 34161 13481 34195 13515
rect 34195 13481 34204 13515
rect 34152 13472 34204 13481
rect 33876 13404 33928 13456
rect 34060 13404 34112 13456
rect 35164 13404 35216 13456
rect 31024 13336 31076 13388
rect 32496 13336 32548 13388
rect 27804 13268 27856 13320
rect 28632 13200 28684 13252
rect 30472 13132 30524 13184
rect 30748 13200 30800 13252
rect 31024 13200 31076 13252
rect 31208 13268 31260 13320
rect 33876 13311 33928 13320
rect 33876 13277 33885 13311
rect 33885 13277 33919 13311
rect 33919 13277 33928 13311
rect 33876 13268 33928 13277
rect 33968 13311 34020 13320
rect 33968 13277 33977 13311
rect 33977 13277 34011 13311
rect 34011 13277 34020 13311
rect 35624 13336 35676 13388
rect 38108 13379 38160 13388
rect 38108 13345 38117 13379
rect 38117 13345 38151 13379
rect 38151 13345 38160 13379
rect 38108 13336 38160 13345
rect 33968 13268 34020 13277
rect 34796 13268 34848 13320
rect 35256 13268 35308 13320
rect 35992 13268 36044 13320
rect 35164 13200 35216 13252
rect 31392 13132 31444 13184
rect 34152 13132 34204 13184
rect 34520 13132 34572 13184
rect 35348 13132 35400 13184
rect 37648 13200 37700 13252
rect 36268 13132 36320 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 16120 12928 16172 12980
rect 18696 12928 18748 12980
rect 19340 12928 19392 12980
rect 20720 12928 20772 12980
rect 26424 12928 26476 12980
rect 34060 12928 34112 12980
rect 36452 12928 36504 12980
rect 37648 12971 37700 12980
rect 37648 12937 37657 12971
rect 37657 12937 37691 12971
rect 37691 12937 37700 12971
rect 37648 12928 37700 12937
rect 13820 12860 13872 12912
rect 17132 12860 17184 12912
rect 19064 12903 19116 12912
rect 19064 12869 19073 12903
rect 19073 12869 19107 12903
rect 19107 12869 19116 12903
rect 19064 12860 19116 12869
rect 19156 12903 19208 12912
rect 19156 12869 19165 12903
rect 19165 12869 19199 12903
rect 19199 12869 19208 12903
rect 19156 12860 19208 12869
rect 2964 12792 3016 12844
rect 4068 12792 4120 12844
rect 15200 12792 15252 12844
rect 16672 12792 16724 12844
rect 16764 12792 16816 12844
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 18696 12792 18748 12844
rect 20996 12903 21048 12912
rect 20996 12869 21005 12903
rect 21005 12869 21039 12903
rect 21039 12869 21048 12903
rect 20996 12860 21048 12869
rect 21180 12903 21232 12912
rect 21180 12869 21189 12903
rect 21189 12869 21223 12903
rect 21223 12869 21232 12903
rect 21180 12860 21232 12869
rect 19432 12823 19439 12844
rect 19439 12823 19473 12844
rect 19473 12823 19484 12844
rect 19432 12792 19484 12823
rect 20628 12792 20680 12844
rect 22192 12860 22244 12912
rect 22928 12860 22980 12912
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 22652 12792 22704 12844
rect 23940 12860 23992 12912
rect 24768 12903 24820 12912
rect 24768 12869 24777 12903
rect 24777 12869 24811 12903
rect 24811 12869 24820 12903
rect 24768 12860 24820 12869
rect 26976 12903 27028 12912
rect 26976 12869 26985 12903
rect 26985 12869 27019 12903
rect 27019 12869 27028 12903
rect 26976 12860 27028 12869
rect 28632 12903 28684 12912
rect 28632 12869 28641 12903
rect 28641 12869 28675 12903
rect 28675 12869 28684 12903
rect 28632 12860 28684 12869
rect 31300 12860 31352 12912
rect 23388 12835 23440 12844
rect 23388 12801 23397 12835
rect 23397 12801 23431 12835
rect 23431 12801 23440 12835
rect 24216 12835 24268 12844
rect 23388 12792 23440 12801
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 25780 12792 25832 12844
rect 18788 12724 18840 12776
rect 20904 12724 20956 12776
rect 21088 12724 21140 12776
rect 22928 12724 22980 12776
rect 25320 12724 25372 12776
rect 25504 12724 25556 12776
rect 26792 12792 26844 12844
rect 29552 12835 29604 12844
rect 29552 12801 29561 12835
rect 29561 12801 29595 12835
rect 29595 12801 29604 12835
rect 29552 12792 29604 12801
rect 29736 12835 29788 12844
rect 29736 12801 29745 12835
rect 29745 12801 29779 12835
rect 29779 12801 29788 12835
rect 29736 12792 29788 12801
rect 29920 12835 29972 12844
rect 29920 12801 29929 12835
rect 29929 12801 29963 12835
rect 29963 12801 29972 12835
rect 29920 12792 29972 12801
rect 30932 12792 30984 12844
rect 31208 12835 31260 12844
rect 31208 12801 31217 12835
rect 31217 12801 31251 12835
rect 31251 12801 31260 12835
rect 31208 12792 31260 12801
rect 29644 12767 29696 12776
rect 29644 12733 29653 12767
rect 29653 12733 29687 12767
rect 29687 12733 29696 12767
rect 29644 12724 29696 12733
rect 31116 12767 31168 12776
rect 31116 12733 31125 12767
rect 31125 12733 31159 12767
rect 31159 12733 31168 12767
rect 31116 12724 31168 12733
rect 32036 12860 32088 12912
rect 32404 12860 32456 12912
rect 33692 12860 33744 12912
rect 34520 12860 34572 12912
rect 35716 12860 35768 12912
rect 33600 12792 33652 12844
rect 35348 12835 35400 12844
rect 19340 12656 19392 12708
rect 19984 12656 20036 12708
rect 25688 12656 25740 12708
rect 30288 12656 30340 12708
rect 30380 12656 30432 12708
rect 32404 12724 32456 12776
rect 33876 12724 33928 12776
rect 34612 12724 34664 12776
rect 35348 12801 35357 12835
rect 35357 12801 35391 12835
rect 35391 12801 35400 12835
rect 35348 12792 35400 12801
rect 35808 12835 35860 12844
rect 35808 12801 35817 12835
rect 35817 12801 35851 12835
rect 35851 12801 35860 12835
rect 35808 12792 35860 12801
rect 36084 12860 36136 12912
rect 36636 12835 36688 12844
rect 36636 12801 36645 12835
rect 36645 12801 36679 12835
rect 36679 12801 36688 12835
rect 36636 12792 36688 12801
rect 37556 12835 37608 12844
rect 37556 12801 37565 12835
rect 37565 12801 37599 12835
rect 37599 12801 37608 12835
rect 37556 12792 37608 12801
rect 36084 12724 36136 12776
rect 36268 12724 36320 12776
rect 32496 12656 32548 12708
rect 1584 12588 1636 12640
rect 14004 12631 14056 12640
rect 14004 12597 14013 12631
rect 14013 12597 14047 12631
rect 14047 12597 14056 12631
rect 14004 12588 14056 12597
rect 23480 12631 23532 12640
rect 23480 12597 23489 12631
rect 23489 12597 23523 12631
rect 23523 12597 23532 12631
rect 23480 12588 23532 12597
rect 24124 12631 24176 12640
rect 24124 12597 24133 12631
rect 24133 12597 24167 12631
rect 24167 12597 24176 12631
rect 24124 12588 24176 12597
rect 25780 12631 25832 12640
rect 25780 12597 25789 12631
rect 25789 12597 25823 12631
rect 25823 12597 25832 12631
rect 25780 12588 25832 12597
rect 25964 12588 26016 12640
rect 27712 12631 27764 12640
rect 27712 12597 27721 12631
rect 27721 12597 27755 12631
rect 27755 12597 27764 12631
rect 27712 12588 27764 12597
rect 29460 12631 29512 12640
rect 29460 12597 29469 12631
rect 29469 12597 29503 12631
rect 29503 12597 29512 12631
rect 29460 12588 29512 12597
rect 31852 12588 31904 12640
rect 32312 12631 32364 12640
rect 32312 12597 32321 12631
rect 32321 12597 32355 12631
rect 32355 12597 32364 12631
rect 32312 12588 32364 12597
rect 33968 12588 34020 12640
rect 34612 12588 34664 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 18328 12384 18380 12436
rect 24216 12384 24268 12436
rect 25596 12384 25648 12436
rect 28816 12427 28868 12436
rect 28816 12393 28825 12427
rect 28825 12393 28859 12427
rect 28859 12393 28868 12427
rect 28816 12384 28868 12393
rect 29736 12384 29788 12436
rect 29920 12384 29972 12436
rect 32312 12384 32364 12436
rect 33600 12384 33652 12436
rect 34428 12384 34480 12436
rect 35624 12384 35676 12436
rect 17040 12316 17092 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 1584 12291 1636 12300
rect 1584 12257 1593 12291
rect 1593 12257 1627 12291
rect 1627 12257 1636 12291
rect 1584 12248 1636 12257
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 16764 12248 16816 12300
rect 17960 12248 18012 12300
rect 18696 12248 18748 12300
rect 22836 12316 22888 12368
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 18052 12180 18104 12232
rect 14004 12112 14056 12164
rect 14372 12044 14424 12096
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 17776 12044 17828 12096
rect 18788 12112 18840 12164
rect 19248 12112 19300 12164
rect 20076 12180 20128 12232
rect 23480 12248 23532 12300
rect 25964 12248 26016 12300
rect 32404 12291 32456 12300
rect 20904 12180 20956 12232
rect 21180 12180 21232 12232
rect 21916 12223 21968 12232
rect 21916 12189 21925 12223
rect 21925 12189 21959 12223
rect 21959 12189 21968 12223
rect 21916 12180 21968 12189
rect 22376 12223 22428 12232
rect 22376 12189 22385 12223
rect 22385 12189 22419 12223
rect 22419 12189 22428 12223
rect 22376 12180 22428 12189
rect 22928 12180 22980 12232
rect 24768 12180 24820 12232
rect 25412 12180 25464 12232
rect 26332 12180 26384 12232
rect 26608 12223 26660 12232
rect 26608 12189 26617 12223
rect 26617 12189 26651 12223
rect 26651 12189 26660 12223
rect 26608 12180 26660 12189
rect 29000 12223 29052 12232
rect 29000 12189 29009 12223
rect 29009 12189 29043 12223
rect 29043 12189 29052 12223
rect 29000 12180 29052 12189
rect 20628 12044 20680 12096
rect 23572 12112 23624 12164
rect 27620 12112 27672 12164
rect 30380 12180 30432 12232
rect 30472 12223 30524 12232
rect 30472 12189 30481 12223
rect 30481 12189 30515 12223
rect 30515 12189 30524 12223
rect 30932 12223 30984 12232
rect 30472 12180 30524 12189
rect 30932 12189 30941 12223
rect 30941 12189 30975 12223
rect 30975 12189 30984 12223
rect 30932 12180 30984 12189
rect 31024 12180 31076 12232
rect 32404 12257 32413 12291
rect 32413 12257 32447 12291
rect 32447 12257 32456 12291
rect 32404 12248 32456 12257
rect 34152 12180 34204 12232
rect 36820 12248 36872 12300
rect 36268 12223 36320 12232
rect 36268 12189 36277 12223
rect 36277 12189 36311 12223
rect 36311 12189 36320 12223
rect 36268 12180 36320 12189
rect 30748 12112 30800 12164
rect 31208 12155 31260 12164
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 29368 12044 29420 12096
rect 31208 12121 31217 12155
rect 31217 12121 31251 12155
rect 31251 12121 31260 12155
rect 31208 12112 31260 12121
rect 31116 12087 31168 12096
rect 31116 12053 31125 12087
rect 31125 12053 31159 12087
rect 31159 12053 31168 12087
rect 32404 12112 32456 12164
rect 37648 12112 37700 12164
rect 38108 12155 38160 12164
rect 38108 12121 38117 12155
rect 38117 12121 38151 12155
rect 38151 12121 38160 12155
rect 38108 12112 38160 12121
rect 31760 12087 31812 12096
rect 31116 12044 31168 12053
rect 31760 12053 31769 12087
rect 31769 12053 31803 12087
rect 31803 12053 31812 12087
rect 31760 12044 31812 12053
rect 32128 12087 32180 12096
rect 32128 12053 32137 12087
rect 32137 12053 32171 12087
rect 32171 12053 32180 12087
rect 32128 12044 32180 12053
rect 32680 12044 32732 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 13084 11840 13136 11892
rect 13912 11840 13964 11892
rect 17316 11840 17368 11892
rect 17500 11840 17552 11892
rect 17960 11840 18012 11892
rect 18236 11840 18288 11892
rect 18604 11883 18656 11892
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 20628 11840 20680 11892
rect 21916 11840 21968 11892
rect 25780 11883 25832 11892
rect 25780 11849 25789 11883
rect 25789 11849 25823 11883
rect 25823 11849 25832 11883
rect 25780 11840 25832 11849
rect 26792 11840 26844 11892
rect 15200 11772 15252 11824
rect 19064 11772 19116 11824
rect 20444 11772 20496 11824
rect 14280 11704 14332 11756
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 16120 11704 16172 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 18696 11747 18748 11756
rect 1584 11679 1636 11688
rect 1584 11645 1593 11679
rect 1593 11645 1627 11679
rect 1627 11645 1636 11679
rect 1584 11636 1636 11645
rect 1952 11636 2004 11688
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 14188 11636 14240 11688
rect 18052 11636 18104 11688
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 19248 11704 19300 11756
rect 19984 11704 20036 11756
rect 24676 11772 24728 11824
rect 26332 11772 26384 11824
rect 30472 11840 30524 11892
rect 30748 11840 30800 11892
rect 31576 11840 31628 11892
rect 32128 11883 32180 11892
rect 32128 11849 32137 11883
rect 32137 11849 32171 11883
rect 32171 11849 32180 11883
rect 32128 11840 32180 11849
rect 36084 11883 36136 11892
rect 36084 11849 36093 11883
rect 36093 11849 36127 11883
rect 36127 11849 36136 11883
rect 36084 11840 36136 11849
rect 37648 11883 37700 11892
rect 37648 11849 37657 11883
rect 37657 11849 37691 11883
rect 37691 11849 37700 11883
rect 37648 11840 37700 11849
rect 29460 11815 29512 11824
rect 29460 11781 29469 11815
rect 29469 11781 29503 11815
rect 29503 11781 29512 11815
rect 29460 11772 29512 11781
rect 29920 11772 29972 11824
rect 32036 11772 32088 11824
rect 32496 11815 32548 11824
rect 32496 11781 32505 11815
rect 32505 11781 32539 11815
rect 32539 11781 32548 11815
rect 32496 11772 32548 11781
rect 34612 11815 34664 11824
rect 34612 11781 34621 11815
rect 34621 11781 34655 11815
rect 34655 11781 34664 11815
rect 34612 11772 34664 11781
rect 35348 11772 35400 11824
rect 19432 11636 19484 11688
rect 21456 11636 21508 11688
rect 31852 11704 31904 11756
rect 32956 11747 33008 11756
rect 32956 11713 32965 11747
rect 32965 11713 32999 11747
rect 32999 11713 33008 11747
rect 32956 11704 33008 11713
rect 36728 11747 36780 11756
rect 36728 11713 36737 11747
rect 36737 11713 36771 11747
rect 36771 11713 36780 11747
rect 37740 11747 37792 11756
rect 36728 11704 36780 11713
rect 37740 11713 37749 11747
rect 37749 11713 37783 11747
rect 37783 11713 37792 11747
rect 37740 11704 37792 11713
rect 16856 11500 16908 11552
rect 18328 11500 18380 11552
rect 18604 11500 18656 11552
rect 20076 11500 20128 11552
rect 20444 11500 20496 11552
rect 20536 11500 20588 11552
rect 22100 11500 22152 11552
rect 22468 11500 22520 11552
rect 22652 11500 22704 11552
rect 24124 11636 24176 11688
rect 25596 11679 25648 11688
rect 25596 11645 25605 11679
rect 25605 11645 25639 11679
rect 25639 11645 25648 11679
rect 25596 11636 25648 11645
rect 26240 11568 26292 11620
rect 26608 11568 26660 11620
rect 27712 11636 27764 11688
rect 28724 11636 28776 11688
rect 24584 11543 24636 11552
rect 24584 11509 24593 11543
rect 24593 11509 24627 11543
rect 24627 11509 24636 11543
rect 24584 11500 24636 11509
rect 28632 11500 28684 11552
rect 31668 11636 31720 11688
rect 31208 11568 31260 11620
rect 30840 11500 30892 11552
rect 31576 11543 31628 11552
rect 31576 11509 31585 11543
rect 31585 11509 31619 11543
rect 31619 11509 31628 11543
rect 31576 11500 31628 11509
rect 33416 11500 33468 11552
rect 35900 11500 35952 11552
rect 36544 11500 36596 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 17316 11296 17368 11348
rect 22468 11296 22520 11348
rect 22928 11296 22980 11348
rect 15936 11160 15988 11212
rect 16396 11160 16448 11212
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2044 11092 2096 11101
rect 2228 11092 2280 11144
rect 14372 11092 14424 11144
rect 15292 11092 15344 11144
rect 17960 11160 18012 11212
rect 18604 11160 18656 11212
rect 17776 11024 17828 11076
rect 18696 11024 18748 11076
rect 20260 11092 20312 11144
rect 20904 11092 20956 11144
rect 21456 11203 21508 11212
rect 21456 11169 21465 11203
rect 21465 11169 21499 11203
rect 21499 11169 21508 11203
rect 21456 11160 21508 11169
rect 20076 11024 20128 11076
rect 21548 11092 21600 11144
rect 24124 11228 24176 11280
rect 23756 11160 23808 11212
rect 24584 11160 24636 11212
rect 24768 11228 24820 11280
rect 25228 11228 25280 11280
rect 26700 11296 26752 11348
rect 27436 11296 27488 11348
rect 29920 11296 29972 11348
rect 30932 11296 30984 11348
rect 34152 11339 34204 11348
rect 34152 11305 34161 11339
rect 34161 11305 34195 11339
rect 34195 11305 34204 11339
rect 34152 11296 34204 11305
rect 35440 11296 35492 11348
rect 29184 11228 29236 11280
rect 34704 11228 34756 11280
rect 36084 11228 36136 11280
rect 36820 11228 36872 11280
rect 25320 11160 25372 11212
rect 26056 11203 26108 11212
rect 26056 11169 26065 11203
rect 26065 11169 26099 11203
rect 26099 11169 26108 11203
rect 26056 11160 26108 11169
rect 18052 10956 18104 11008
rect 20812 10956 20864 11008
rect 22928 11135 22980 11144
rect 22928 11101 22937 11135
rect 22937 11101 22971 11135
rect 22971 11101 22980 11135
rect 23572 11135 23624 11144
rect 22928 11092 22980 11101
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 24032 11092 24084 11144
rect 24308 11092 24360 11144
rect 25964 11135 26016 11144
rect 25964 11101 25973 11135
rect 25973 11101 26007 11135
rect 26007 11101 26016 11135
rect 25964 11092 26016 11101
rect 22192 10956 22244 11008
rect 23848 11024 23900 11076
rect 24952 11024 25004 11076
rect 26700 11092 26752 11144
rect 27252 11160 27304 11212
rect 29368 11160 29420 11212
rect 31668 11160 31720 11212
rect 32680 11203 32732 11212
rect 32680 11169 32689 11203
rect 32689 11169 32723 11203
rect 32723 11169 32732 11203
rect 32680 11160 32732 11169
rect 35440 11160 35492 11212
rect 27068 11092 27120 11144
rect 27804 11092 27856 11144
rect 30380 11092 30432 11144
rect 36084 11092 36136 11144
rect 23388 10956 23440 11008
rect 23664 10956 23716 11008
rect 24308 10956 24360 11008
rect 25412 10956 25464 11008
rect 30932 11024 30984 11076
rect 31576 11024 31628 11076
rect 35624 11024 35676 11076
rect 36636 11024 36688 11076
rect 38200 11024 38252 11076
rect 27252 10956 27304 11008
rect 27896 10956 27948 11008
rect 31024 10956 31076 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 14280 10752 14332 10804
rect 15292 10752 15344 10804
rect 16396 10752 16448 10804
rect 18052 10752 18104 10804
rect 17132 10727 17184 10736
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 17776 10727 17828 10736
rect 17776 10693 17785 10727
rect 17785 10693 17819 10727
rect 17819 10693 17828 10727
rect 17776 10684 17828 10693
rect 18144 10727 18196 10736
rect 18144 10693 18153 10727
rect 18153 10693 18187 10727
rect 18187 10693 18196 10727
rect 18144 10684 18196 10693
rect 18696 10752 18748 10804
rect 22284 10752 22336 10804
rect 22744 10752 22796 10804
rect 23204 10684 23256 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 15200 10616 15252 10668
rect 15384 10616 15436 10668
rect 16672 10616 16724 10668
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 15844 10591 15896 10600
rect 15844 10557 15853 10591
rect 15853 10557 15887 10591
rect 15887 10557 15896 10591
rect 15844 10548 15896 10557
rect 17684 10548 17736 10600
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 22100 10616 22152 10668
rect 23940 10684 23992 10736
rect 24124 10727 24176 10736
rect 24124 10693 24133 10727
rect 24133 10693 24167 10727
rect 24167 10693 24176 10727
rect 24124 10684 24176 10693
rect 24308 10727 24360 10736
rect 24308 10693 24333 10727
rect 24333 10693 24360 10727
rect 25964 10752 26016 10804
rect 27620 10752 27672 10804
rect 29184 10795 29236 10804
rect 29184 10761 29193 10795
rect 29193 10761 29227 10795
rect 29227 10761 29236 10795
rect 29184 10752 29236 10761
rect 30380 10752 30432 10804
rect 24308 10684 24360 10693
rect 25412 10684 25464 10736
rect 26976 10684 27028 10736
rect 23388 10659 23440 10668
rect 23388 10625 23397 10659
rect 23397 10625 23431 10659
rect 23431 10625 23440 10659
rect 23388 10616 23440 10625
rect 23664 10616 23716 10668
rect 24584 10616 24636 10668
rect 25228 10659 25280 10668
rect 25228 10625 25237 10659
rect 25237 10625 25271 10659
rect 25271 10625 25280 10659
rect 25228 10616 25280 10625
rect 25596 10616 25648 10668
rect 28172 10684 28224 10736
rect 29276 10684 29328 10736
rect 29828 10684 29880 10736
rect 27252 10659 27304 10668
rect 27252 10625 27261 10659
rect 27261 10625 27295 10659
rect 27295 10625 27304 10659
rect 27252 10616 27304 10625
rect 28080 10616 28132 10668
rect 16856 10480 16908 10532
rect 19892 10548 19944 10600
rect 20628 10548 20680 10600
rect 20996 10591 21048 10600
rect 20996 10557 21005 10591
rect 21005 10557 21039 10591
rect 21039 10557 21048 10591
rect 20996 10548 21048 10557
rect 22008 10548 22060 10600
rect 24676 10548 24728 10600
rect 15568 10412 15620 10464
rect 16764 10412 16816 10464
rect 19432 10412 19484 10464
rect 19708 10412 19760 10464
rect 20536 10412 20588 10464
rect 20904 10480 20956 10532
rect 23388 10480 23440 10532
rect 24124 10480 24176 10532
rect 24952 10523 25004 10532
rect 24952 10489 24961 10523
rect 24961 10489 24995 10523
rect 24995 10489 25004 10523
rect 24952 10480 25004 10489
rect 26148 10480 26200 10532
rect 28172 10548 28224 10600
rect 28632 10616 28684 10668
rect 30840 10684 30892 10736
rect 31668 10752 31720 10804
rect 33876 10795 33928 10804
rect 33876 10761 33885 10795
rect 33885 10761 33919 10795
rect 33919 10761 33928 10795
rect 33876 10752 33928 10761
rect 31392 10684 31444 10736
rect 33416 10684 33468 10736
rect 36544 10727 36596 10736
rect 36544 10693 36553 10727
rect 36553 10693 36587 10727
rect 36587 10693 36596 10727
rect 36544 10684 36596 10693
rect 38568 10616 38620 10668
rect 30196 10548 30248 10600
rect 31668 10548 31720 10600
rect 35808 10591 35860 10600
rect 35808 10557 35817 10591
rect 35817 10557 35851 10591
rect 35851 10557 35860 10591
rect 35808 10548 35860 10557
rect 36728 10591 36780 10600
rect 36728 10557 36737 10591
rect 36737 10557 36771 10591
rect 36771 10557 36780 10591
rect 36728 10548 36780 10557
rect 32128 10480 32180 10532
rect 21548 10412 21600 10464
rect 22744 10412 22796 10464
rect 25228 10412 25280 10464
rect 26240 10412 26292 10464
rect 29368 10455 29420 10464
rect 29368 10421 29377 10455
rect 29377 10421 29411 10455
rect 29411 10421 29420 10455
rect 29368 10412 29420 10421
rect 36452 10412 36504 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 17592 10208 17644 10260
rect 16856 10140 16908 10192
rect 18052 10208 18104 10260
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 20996 10208 21048 10260
rect 22652 10208 22704 10260
rect 23572 10251 23624 10260
rect 23572 10217 23581 10251
rect 23581 10217 23615 10251
rect 23615 10217 23624 10251
rect 23572 10208 23624 10217
rect 15200 10004 15252 10056
rect 15384 10004 15436 10056
rect 16580 10004 16632 10056
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 20076 10140 20128 10192
rect 22100 10140 22152 10192
rect 18788 10072 18840 10124
rect 17316 10004 17368 10013
rect 18972 10004 19024 10056
rect 22008 10072 22060 10124
rect 22744 10115 22796 10124
rect 22744 10081 22753 10115
rect 22753 10081 22787 10115
rect 22787 10081 22796 10115
rect 22744 10072 22796 10081
rect 18328 9936 18380 9988
rect 18880 9936 18932 9988
rect 19156 9936 19208 9988
rect 23480 10004 23532 10056
rect 27804 10251 27856 10260
rect 27804 10217 27813 10251
rect 27813 10217 27847 10251
rect 27847 10217 27856 10251
rect 27804 10208 27856 10217
rect 27896 10208 27948 10260
rect 30196 10208 30248 10260
rect 30932 10251 30984 10260
rect 30932 10217 30941 10251
rect 30941 10217 30975 10251
rect 30975 10217 30984 10251
rect 30932 10208 30984 10217
rect 31668 10251 31720 10260
rect 31668 10217 31677 10251
rect 31677 10217 31711 10251
rect 31711 10217 31720 10251
rect 31668 10208 31720 10217
rect 32128 10208 32180 10260
rect 35348 10208 35400 10260
rect 35624 10251 35676 10260
rect 35624 10217 35633 10251
rect 35633 10217 35667 10251
rect 35667 10217 35676 10251
rect 35624 10208 35676 10217
rect 26332 10140 26384 10192
rect 29000 10140 29052 10192
rect 26240 10072 26292 10124
rect 27528 10072 27580 10124
rect 28172 10115 28224 10124
rect 28172 10081 28181 10115
rect 28181 10081 28215 10115
rect 28215 10081 28224 10115
rect 28172 10072 28224 10081
rect 20444 9979 20496 9988
rect 20444 9945 20453 9979
rect 20453 9945 20487 9979
rect 20487 9945 20496 9979
rect 20444 9936 20496 9945
rect 22192 9979 22244 9988
rect 22192 9945 22201 9979
rect 22201 9945 22235 9979
rect 22235 9945 22244 9979
rect 22192 9936 22244 9945
rect 27896 10004 27948 10056
rect 28080 10047 28132 10056
rect 28080 10013 28089 10047
rect 28089 10013 28123 10047
rect 28123 10013 28132 10047
rect 28080 10004 28132 10013
rect 28264 10004 28316 10056
rect 29644 10004 29696 10056
rect 29828 10047 29880 10056
rect 29828 10013 29837 10047
rect 29837 10013 29871 10047
rect 29871 10013 29880 10047
rect 29828 10004 29880 10013
rect 30380 10004 30432 10056
rect 36452 10115 36504 10124
rect 36452 10081 36461 10115
rect 36461 10081 36495 10115
rect 36495 10081 36504 10115
rect 36452 10072 36504 10081
rect 38108 10115 38160 10124
rect 38108 10081 38117 10115
rect 38117 10081 38151 10115
rect 38151 10081 38160 10115
rect 38108 10072 38160 10081
rect 31760 10004 31812 10056
rect 25228 9979 25280 9988
rect 25228 9945 25237 9979
rect 25237 9945 25271 9979
rect 25271 9945 25280 9979
rect 25228 9936 25280 9945
rect 28540 9936 28592 9988
rect 29000 9979 29052 9988
rect 29000 9945 29009 9979
rect 29009 9945 29043 9979
rect 29043 9945 29052 9979
rect 29000 9936 29052 9945
rect 31024 9936 31076 9988
rect 32956 10004 33008 10056
rect 14096 9868 14148 9920
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 19248 9868 19300 9920
rect 22652 9911 22704 9920
rect 22652 9877 22661 9911
rect 22661 9877 22695 9911
rect 22695 9877 22704 9911
rect 22652 9868 22704 9877
rect 23388 9911 23440 9920
rect 23388 9877 23397 9911
rect 23397 9877 23431 9911
rect 23431 9877 23440 9911
rect 23388 9868 23440 9877
rect 23848 9868 23900 9920
rect 26700 9911 26752 9920
rect 26700 9877 26709 9911
rect 26709 9877 26743 9911
rect 26743 9877 26752 9911
rect 26700 9868 26752 9877
rect 27896 9868 27948 9920
rect 30380 9868 30432 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 18052 9707 18104 9716
rect 18052 9673 18061 9707
rect 18061 9673 18095 9707
rect 18095 9673 18104 9707
rect 18052 9664 18104 9673
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 20812 9707 20864 9716
rect 14096 9596 14148 9648
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 16856 9596 16908 9648
rect 16948 9596 17000 9648
rect 17960 9596 18012 9648
rect 18696 9596 18748 9648
rect 20812 9673 20821 9707
rect 20821 9673 20855 9707
rect 20855 9673 20864 9707
rect 20812 9664 20864 9673
rect 20904 9664 20956 9716
rect 13452 9460 13504 9512
rect 19248 9596 19300 9648
rect 25228 9664 25280 9716
rect 17408 9528 17460 9580
rect 18880 9571 18932 9580
rect 18880 9537 18889 9571
rect 18889 9537 18923 9571
rect 18923 9537 18932 9571
rect 18880 9528 18932 9537
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 19156 9528 19208 9580
rect 15476 9392 15528 9444
rect 16580 9460 16632 9512
rect 17224 9460 17276 9512
rect 18052 9460 18104 9512
rect 19892 9528 19944 9580
rect 20076 9528 20128 9580
rect 21456 9528 21508 9580
rect 22560 9596 22612 9648
rect 23388 9596 23440 9648
rect 22468 9528 22520 9580
rect 25688 9596 25740 9648
rect 25964 9596 26016 9648
rect 28264 9664 28316 9716
rect 30196 9664 30248 9716
rect 27528 9639 27580 9648
rect 18604 9392 18656 9444
rect 20904 9460 20956 9512
rect 21180 9503 21232 9512
rect 21180 9469 21189 9503
rect 21189 9469 21223 9503
rect 21223 9469 21232 9503
rect 21180 9460 21232 9469
rect 22100 9460 22152 9512
rect 23480 9460 23532 9512
rect 1400 9324 1452 9376
rect 4068 9324 4120 9376
rect 16580 9324 16632 9376
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 19340 9324 19392 9376
rect 19984 9367 20036 9376
rect 19984 9333 19993 9367
rect 19993 9333 20027 9367
rect 20027 9333 20036 9367
rect 19984 9324 20036 9333
rect 20904 9324 20956 9376
rect 21548 9324 21600 9376
rect 22744 9324 22796 9376
rect 23756 9392 23808 9444
rect 24124 9571 24176 9580
rect 24124 9537 24133 9571
rect 24133 9537 24167 9571
rect 24167 9537 24176 9571
rect 24124 9528 24176 9537
rect 25320 9528 25372 9580
rect 25872 9528 25924 9580
rect 26424 9528 26476 9580
rect 27160 9528 27212 9580
rect 27528 9605 27537 9639
rect 27537 9605 27571 9639
rect 27571 9605 27580 9639
rect 27528 9596 27580 9605
rect 27436 9571 27488 9580
rect 27436 9537 27453 9571
rect 27453 9537 27488 9571
rect 27436 9528 27488 9537
rect 24676 9460 24728 9512
rect 25964 9503 26016 9512
rect 24124 9392 24176 9444
rect 23664 9367 23716 9376
rect 23664 9333 23673 9367
rect 23673 9333 23707 9367
rect 23707 9333 23716 9367
rect 25044 9367 25096 9376
rect 23664 9324 23716 9333
rect 25044 9333 25053 9367
rect 25053 9333 25087 9367
rect 25087 9333 25096 9367
rect 25044 9324 25096 9333
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 26148 9503 26200 9512
rect 26148 9469 26157 9503
rect 26157 9469 26191 9503
rect 26191 9469 26200 9503
rect 26148 9460 26200 9469
rect 26240 9503 26292 9512
rect 26240 9469 26249 9503
rect 26249 9469 26283 9503
rect 26283 9469 26292 9503
rect 26240 9460 26292 9469
rect 26516 9460 26568 9512
rect 30472 9596 30524 9648
rect 36636 9639 36688 9648
rect 36636 9605 36645 9639
rect 36645 9605 36679 9639
rect 36679 9605 36688 9639
rect 36636 9596 36688 9605
rect 30012 9528 30064 9580
rect 31024 9571 31076 9580
rect 31024 9537 31033 9571
rect 31033 9537 31067 9571
rect 31067 9537 31076 9571
rect 31024 9528 31076 9537
rect 35992 9528 36044 9580
rect 37004 9528 37056 9580
rect 38384 9528 38436 9580
rect 27896 9460 27948 9512
rect 28632 9503 28684 9512
rect 28632 9469 28641 9503
rect 28641 9469 28675 9503
rect 28675 9469 28684 9503
rect 28632 9460 28684 9469
rect 36176 9460 36228 9512
rect 36268 9392 36320 9444
rect 26976 9324 27028 9376
rect 37924 9324 37976 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 15476 9120 15528 9172
rect 15844 9120 15896 9172
rect 18052 9120 18104 9172
rect 17040 9052 17092 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 15936 8984 15988 9036
rect 17500 8984 17552 9036
rect 17868 9052 17920 9104
rect 19248 9120 19300 9172
rect 20904 9120 20956 9172
rect 19432 9052 19484 9104
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 5816 8916 5868 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 1952 8848 2004 8900
rect 14832 8848 14884 8900
rect 17224 8959 17276 8968
rect 17224 8925 17233 8959
rect 17233 8925 17267 8959
rect 17267 8925 17276 8959
rect 17592 8959 17644 8968
rect 17224 8916 17276 8925
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 17960 8916 18012 8968
rect 18144 8916 18196 8968
rect 16856 8848 16908 8900
rect 4344 8780 4396 8832
rect 17132 8780 17184 8832
rect 17868 8848 17920 8900
rect 18328 8891 18380 8900
rect 18328 8857 18337 8891
rect 18337 8857 18371 8891
rect 18371 8857 18380 8891
rect 18328 8848 18380 8857
rect 18788 8916 18840 8968
rect 19984 8916 20036 8968
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 22100 9120 22152 9172
rect 22008 9052 22060 9104
rect 22744 9163 22796 9172
rect 22744 9129 22753 9163
rect 22753 9129 22787 9163
rect 22787 9129 22796 9163
rect 22744 9120 22796 9129
rect 25044 9120 25096 9172
rect 30012 9120 30064 9172
rect 35440 9163 35492 9172
rect 35440 9129 35449 9163
rect 35449 9129 35483 9163
rect 35483 9129 35492 9163
rect 35440 9120 35492 9129
rect 22928 9052 22980 9104
rect 23112 9052 23164 9104
rect 24676 9052 24728 9104
rect 25780 9052 25832 9104
rect 26056 9052 26108 9104
rect 27436 9052 27488 9104
rect 21272 8984 21324 8993
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 22192 8959 22244 8968
rect 21456 8916 21508 8925
rect 18880 8780 18932 8832
rect 20628 8848 20680 8900
rect 22192 8925 22201 8959
rect 22201 8925 22235 8959
rect 22235 8925 22244 8959
rect 22192 8916 22244 8925
rect 22284 8916 22336 8968
rect 22836 8916 22888 8968
rect 24492 8984 24544 9036
rect 25044 8984 25096 9036
rect 25596 8984 25648 9036
rect 26424 8984 26476 9036
rect 28540 9052 28592 9104
rect 37188 9027 37240 9036
rect 20076 8780 20128 8832
rect 22468 8848 22520 8900
rect 25136 8916 25188 8968
rect 26056 8959 26108 8968
rect 26056 8925 26065 8959
rect 26065 8925 26099 8959
rect 26099 8925 26108 8959
rect 26056 8916 26108 8925
rect 24768 8891 24820 8900
rect 24768 8857 24777 8891
rect 24777 8857 24811 8891
rect 24811 8857 24820 8891
rect 24768 8848 24820 8857
rect 22744 8780 22796 8832
rect 24400 8823 24452 8832
rect 24400 8789 24409 8823
rect 24409 8789 24443 8823
rect 24443 8789 24452 8823
rect 24400 8780 24452 8789
rect 24676 8823 24728 8832
rect 24676 8789 24685 8823
rect 24685 8789 24719 8823
rect 24719 8789 24728 8823
rect 27804 8916 27856 8968
rect 28264 8916 28316 8968
rect 37188 8993 37197 9027
rect 37197 8993 37231 9027
rect 37231 8993 37240 9027
rect 37188 8984 37240 8993
rect 37924 9027 37976 9036
rect 37924 8993 37933 9027
rect 37933 8993 37967 9027
rect 37967 8993 37976 9027
rect 37924 8984 37976 8993
rect 29644 8916 29696 8968
rect 30196 8916 30248 8968
rect 30380 8916 30432 8968
rect 38108 8959 38160 8968
rect 38108 8925 38117 8959
rect 38117 8925 38151 8959
rect 38151 8925 38160 8959
rect 38108 8916 38160 8925
rect 26884 8891 26936 8900
rect 26884 8857 26893 8891
rect 26893 8857 26927 8891
rect 26927 8857 26936 8891
rect 26884 8848 26936 8857
rect 24676 8780 24728 8789
rect 26240 8780 26292 8832
rect 26424 8823 26476 8832
rect 26424 8789 26433 8823
rect 26433 8789 26467 8823
rect 26467 8789 26476 8823
rect 26424 8780 26476 8789
rect 26792 8780 26844 8832
rect 27436 8891 27488 8900
rect 27436 8857 27445 8891
rect 27445 8857 27479 8891
rect 27479 8857 27488 8891
rect 27436 8848 27488 8857
rect 27988 8848 28040 8900
rect 27620 8780 27672 8832
rect 28080 8780 28132 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 13544 8576 13596 8628
rect 16672 8619 16724 8628
rect 16672 8585 16681 8619
rect 16681 8585 16715 8619
rect 16715 8585 16724 8619
rect 16672 8576 16724 8585
rect 17408 8576 17460 8628
rect 18236 8576 18288 8628
rect 20352 8576 20404 8628
rect 22836 8619 22888 8628
rect 4344 8551 4396 8560
rect 4344 8517 4353 8551
rect 4353 8517 4387 8551
rect 4387 8517 4396 8551
rect 4344 8508 4396 8517
rect 2136 8440 2188 8492
rect 7932 8440 7984 8492
rect 9956 8440 10008 8492
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17500 8440 17552 8492
rect 18788 8551 18840 8560
rect 18788 8517 18815 8551
rect 18815 8517 18840 8551
rect 18788 8508 18840 8517
rect 19064 8508 19116 8560
rect 19432 8508 19484 8560
rect 22836 8585 22845 8619
rect 22845 8585 22879 8619
rect 22879 8585 22888 8619
rect 22836 8576 22888 8585
rect 23940 8619 23992 8628
rect 23940 8585 23949 8619
rect 23949 8585 23983 8619
rect 23983 8585 23992 8619
rect 23940 8576 23992 8585
rect 24676 8576 24728 8628
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 25136 8576 25188 8628
rect 26884 8576 26936 8628
rect 27804 8576 27856 8628
rect 29644 8576 29696 8628
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 19340 8440 19392 8492
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 4068 8372 4120 8424
rect 15384 8372 15436 8424
rect 15660 8372 15712 8424
rect 5632 8304 5684 8356
rect 16948 8304 17000 8356
rect 20076 8440 20128 8492
rect 20536 8440 20588 8492
rect 21180 8440 21232 8492
rect 23112 8508 23164 8560
rect 23204 8508 23256 8560
rect 25044 8551 25096 8560
rect 25044 8517 25053 8551
rect 25053 8517 25087 8551
rect 25087 8517 25096 8551
rect 25044 8508 25096 8517
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 22836 8440 22888 8492
rect 23296 8440 23348 8492
rect 24768 8483 24820 8492
rect 23848 8372 23900 8424
rect 24768 8449 24777 8483
rect 24777 8449 24811 8483
rect 24811 8449 24820 8483
rect 24768 8440 24820 8449
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 26424 8508 26476 8560
rect 30932 8508 30984 8560
rect 26332 8440 26384 8492
rect 27620 8440 27672 8492
rect 36728 8483 36780 8492
rect 36728 8449 36737 8483
rect 36737 8449 36771 8483
rect 36771 8449 36780 8483
rect 36728 8440 36780 8449
rect 38108 8440 38160 8492
rect 25228 8372 25280 8424
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 18052 8304 18104 8356
rect 18236 8304 18288 8356
rect 20628 8304 20680 8356
rect 23756 8304 23808 8356
rect 24308 8304 24360 8356
rect 25872 8304 25924 8356
rect 27804 8372 27856 8424
rect 28724 8415 28776 8424
rect 28724 8381 28733 8415
rect 28733 8381 28767 8415
rect 28767 8381 28776 8415
rect 28724 8372 28776 8381
rect 27620 8304 27672 8356
rect 22376 8236 22428 8288
rect 23480 8236 23532 8288
rect 24032 8236 24084 8288
rect 24768 8236 24820 8288
rect 25320 8236 25372 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 15200 8032 15252 8084
rect 18144 8032 18196 8084
rect 18512 8032 18564 8084
rect 2136 7964 2188 8016
rect 3976 7939 4028 7948
rect 3976 7905 3985 7939
rect 3985 7905 4019 7939
rect 4019 7905 4028 7939
rect 3976 7896 4028 7905
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 18788 7964 18840 8016
rect 21456 7964 21508 8016
rect 22652 8032 22704 8084
rect 25044 8032 25096 8084
rect 26056 8032 26108 8084
rect 30932 8075 30984 8084
rect 30932 8041 30941 8075
rect 30941 8041 30975 8075
rect 30975 8041 30984 8075
rect 30932 8032 30984 8041
rect 38016 8032 38068 8084
rect 22100 7964 22152 8016
rect 25504 7964 25556 8016
rect 25872 7964 25924 8016
rect 22192 7896 22244 7948
rect 26424 7964 26476 8016
rect 27528 7964 27580 8016
rect 27804 7964 27856 8016
rect 26332 7896 26384 7948
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 15752 7828 15804 7880
rect 16396 7871 16448 7880
rect 15752 7692 15804 7744
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 18696 7828 18748 7880
rect 17868 7803 17920 7812
rect 17868 7769 17877 7803
rect 17877 7769 17911 7803
rect 17911 7769 17920 7803
rect 17868 7760 17920 7769
rect 17960 7760 18012 7812
rect 19340 7760 19392 7812
rect 18236 7692 18288 7744
rect 20812 7828 20864 7880
rect 22376 7871 22428 7880
rect 20720 7760 20772 7812
rect 20996 7760 21048 7812
rect 22376 7837 22385 7871
rect 22385 7837 22419 7871
rect 22419 7837 22428 7871
rect 22376 7828 22428 7837
rect 24400 7828 24452 7880
rect 22928 7803 22980 7812
rect 22928 7769 22937 7803
rect 22937 7769 22971 7803
rect 22971 7769 22980 7803
rect 22928 7760 22980 7769
rect 23388 7760 23440 7812
rect 23480 7803 23532 7812
rect 23480 7769 23489 7803
rect 23489 7769 23523 7803
rect 23523 7769 23532 7803
rect 23480 7760 23532 7769
rect 25136 7828 25188 7880
rect 25688 7828 25740 7880
rect 25044 7803 25096 7812
rect 25044 7769 25053 7803
rect 25053 7769 25087 7803
rect 25087 7769 25096 7803
rect 25320 7803 25372 7812
rect 25044 7760 25096 7769
rect 25320 7769 25329 7803
rect 25329 7769 25363 7803
rect 25363 7769 25372 7803
rect 25320 7760 25372 7769
rect 23848 7692 23900 7744
rect 24768 7735 24820 7744
rect 24768 7701 24777 7735
rect 24777 7701 24811 7735
rect 24811 7701 24820 7735
rect 24768 7692 24820 7701
rect 25228 7692 25280 7744
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 26792 7760 26844 7812
rect 26976 7828 27028 7880
rect 27160 7871 27212 7880
rect 27160 7837 27169 7871
rect 27169 7837 27203 7871
rect 27203 7837 27212 7871
rect 27160 7828 27212 7837
rect 27252 7803 27304 7812
rect 27252 7769 27261 7803
rect 27261 7769 27295 7803
rect 27295 7769 27304 7803
rect 27252 7760 27304 7769
rect 27528 7828 27580 7880
rect 27804 7760 27856 7812
rect 27896 7760 27948 7812
rect 28264 7828 28316 7880
rect 30196 7871 30248 7880
rect 30196 7837 30205 7871
rect 30205 7837 30239 7871
rect 30239 7837 30248 7871
rect 30196 7828 30248 7837
rect 30380 7828 30432 7880
rect 35624 7871 35676 7880
rect 35624 7837 35633 7871
rect 35633 7837 35667 7871
rect 35667 7837 35676 7871
rect 35624 7828 35676 7837
rect 28448 7760 28500 7812
rect 38660 7760 38712 7812
rect 27620 7692 27672 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 16396 7488 16448 7540
rect 18420 7488 18472 7540
rect 18880 7488 18932 7540
rect 20076 7531 20128 7540
rect 20076 7497 20085 7531
rect 20085 7497 20119 7531
rect 20119 7497 20128 7531
rect 20076 7488 20128 7497
rect 22192 7531 22244 7540
rect 22192 7497 22201 7531
rect 22201 7497 22235 7531
rect 22235 7497 22244 7531
rect 22192 7488 22244 7497
rect 23572 7488 23624 7540
rect 25044 7488 25096 7540
rect 26424 7488 26476 7540
rect 16948 7420 17000 7472
rect 17684 7420 17736 7472
rect 18512 7420 18564 7472
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 18972 7352 19024 7404
rect 19432 7395 19484 7404
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 16856 7216 16908 7268
rect 17040 7284 17092 7336
rect 18512 7284 18564 7336
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 20720 7420 20772 7472
rect 20904 7463 20956 7472
rect 20904 7429 20913 7463
rect 20913 7429 20947 7463
rect 20947 7429 20956 7463
rect 20904 7420 20956 7429
rect 21456 7420 21508 7472
rect 22376 7420 22428 7472
rect 27252 7488 27304 7540
rect 19524 7352 19576 7361
rect 20168 7395 20220 7404
rect 20168 7361 20177 7395
rect 20177 7361 20211 7395
rect 20211 7361 20220 7395
rect 20168 7352 20220 7361
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 22008 7395 22060 7404
rect 20352 7284 20404 7336
rect 17684 7216 17736 7268
rect 19340 7216 19392 7268
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 23020 7352 23072 7404
rect 23204 7395 23256 7404
rect 23204 7361 23213 7395
rect 23213 7361 23247 7395
rect 23247 7361 23256 7395
rect 23204 7352 23256 7361
rect 23296 7352 23348 7404
rect 24492 7352 24544 7404
rect 24860 7352 24912 7404
rect 25136 7395 25188 7404
rect 25136 7361 25145 7395
rect 25145 7361 25179 7395
rect 25179 7361 25188 7395
rect 25136 7352 25188 7361
rect 25780 7352 25832 7404
rect 26148 7395 26200 7404
rect 26148 7361 26157 7395
rect 26157 7361 26191 7395
rect 26191 7361 26200 7395
rect 26148 7352 26200 7361
rect 26332 7352 26384 7404
rect 27068 7352 27120 7404
rect 27344 7352 27396 7404
rect 28448 7488 28500 7540
rect 27804 7420 27856 7472
rect 29644 7352 29696 7404
rect 35624 7395 35676 7404
rect 35624 7361 35633 7395
rect 35633 7361 35667 7395
rect 35667 7361 35676 7395
rect 35624 7352 35676 7361
rect 22100 7284 22152 7336
rect 22744 7327 22796 7336
rect 22744 7293 22753 7327
rect 22753 7293 22787 7327
rect 22787 7293 22796 7327
rect 22744 7284 22796 7293
rect 24124 7284 24176 7336
rect 27436 7284 27488 7336
rect 27712 7284 27764 7336
rect 28264 7327 28316 7336
rect 28264 7293 28273 7327
rect 28273 7293 28307 7327
rect 28307 7293 28316 7327
rect 28264 7284 28316 7293
rect 22928 7216 22980 7268
rect 23848 7259 23900 7268
rect 23848 7225 23857 7259
rect 23857 7225 23891 7259
rect 23891 7225 23900 7259
rect 23848 7216 23900 7225
rect 25320 7216 25372 7268
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 18420 7148 18472 7200
rect 18512 7148 18564 7200
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 23204 7191 23256 7200
rect 23204 7157 23213 7191
rect 23213 7157 23247 7191
rect 23247 7157 23256 7191
rect 23204 7148 23256 7157
rect 24768 7148 24820 7200
rect 26240 7148 26292 7200
rect 26976 7191 27028 7200
rect 26976 7157 26985 7191
rect 26985 7157 27019 7191
rect 27019 7157 27028 7191
rect 26976 7148 27028 7157
rect 29000 7148 29052 7200
rect 36268 7148 36320 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1952 6944 2004 6996
rect 22744 6944 22796 6996
rect 26792 6944 26844 6996
rect 27896 6944 27948 6996
rect 15844 6808 15896 6860
rect 16672 6808 16724 6860
rect 17040 6808 17092 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 20628 6808 20680 6860
rect 21272 6808 21324 6860
rect 23204 6808 23256 6860
rect 25504 6851 25556 6860
rect 25504 6817 25513 6851
rect 25513 6817 25547 6851
rect 25547 6817 25556 6851
rect 25504 6808 25556 6817
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 16948 6783 17000 6792
rect 16948 6749 16957 6783
rect 16957 6749 16991 6783
rect 16991 6749 17000 6783
rect 16948 6740 17000 6749
rect 18420 6740 18472 6792
rect 20904 6783 20956 6792
rect 5632 6672 5684 6724
rect 14832 6715 14884 6724
rect 14832 6681 14841 6715
rect 14841 6681 14875 6715
rect 14875 6681 14884 6715
rect 14832 6672 14884 6681
rect 15476 6672 15528 6724
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 21088 6783 21140 6792
rect 21088 6749 21097 6783
rect 21097 6749 21131 6783
rect 21131 6749 21140 6783
rect 21088 6740 21140 6749
rect 21456 6740 21508 6792
rect 22008 6740 22060 6792
rect 22192 6740 22244 6792
rect 23112 6740 23164 6792
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 24676 6740 24728 6792
rect 25044 6740 25096 6792
rect 25228 6740 25280 6792
rect 26332 6783 26384 6792
rect 26332 6749 26341 6783
rect 26341 6749 26375 6783
rect 26375 6749 26384 6783
rect 26332 6740 26384 6749
rect 29000 6808 29052 6860
rect 29644 6851 29696 6860
rect 29644 6817 29653 6851
rect 29653 6817 29687 6851
rect 29687 6817 29696 6851
rect 29644 6808 29696 6817
rect 36268 6851 36320 6860
rect 36268 6817 36277 6851
rect 36277 6817 36311 6851
rect 36311 6817 36320 6851
rect 36268 6808 36320 6817
rect 37188 6851 37240 6860
rect 37188 6817 37197 6851
rect 37197 6817 37231 6851
rect 37231 6817 37240 6851
rect 37188 6808 37240 6817
rect 26976 6783 27028 6792
rect 26976 6749 26985 6783
rect 26985 6749 27019 6783
rect 27019 6749 27028 6783
rect 26976 6740 27028 6749
rect 30380 6740 30432 6792
rect 19984 6672 20036 6724
rect 20996 6715 21048 6724
rect 20996 6681 21005 6715
rect 21005 6681 21039 6715
rect 21039 6681 21048 6715
rect 20996 6672 21048 6681
rect 21180 6715 21232 6724
rect 21180 6681 21215 6715
rect 21215 6681 21232 6715
rect 23296 6715 23348 6724
rect 21180 6672 21232 6681
rect 23296 6681 23305 6715
rect 23305 6681 23339 6715
rect 23339 6681 23348 6715
rect 23296 6672 23348 6681
rect 36452 6715 36504 6724
rect 36452 6681 36461 6715
rect 36461 6681 36495 6715
rect 36495 6681 36504 6715
rect 36452 6672 36504 6681
rect 1860 6604 1912 6656
rect 16764 6647 16816 6656
rect 16764 6613 16773 6647
rect 16773 6613 16807 6647
rect 16807 6613 16816 6647
rect 16764 6604 16816 6613
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 18788 6604 18840 6656
rect 20628 6604 20680 6656
rect 22468 6604 22520 6656
rect 23112 6604 23164 6656
rect 25228 6604 25280 6656
rect 28540 6604 28592 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 14832 6400 14884 6452
rect 17040 6443 17092 6452
rect 17040 6409 17065 6443
rect 17065 6409 17092 6443
rect 17040 6400 17092 6409
rect 17960 6400 18012 6452
rect 20996 6443 21048 6452
rect 1860 6375 1912 6384
rect 1860 6341 1869 6375
rect 1869 6341 1903 6375
rect 1903 6341 1912 6375
rect 1860 6332 1912 6341
rect 16856 6375 16908 6384
rect 16856 6341 16865 6375
rect 16865 6341 16899 6375
rect 16899 6341 16908 6375
rect 16856 6332 16908 6341
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 15384 6264 15436 6316
rect 17684 6307 17736 6316
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 17684 6273 17693 6307
rect 17693 6273 17727 6307
rect 17727 6273 17736 6307
rect 17684 6264 17736 6273
rect 18144 6332 18196 6384
rect 18788 6332 18840 6384
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 19984 6332 20036 6384
rect 20352 6332 20404 6384
rect 20904 6332 20956 6384
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 18512 6264 18564 6316
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 16672 6060 16724 6112
rect 18420 6128 18472 6180
rect 18604 6128 18656 6180
rect 20444 6196 20496 6248
rect 21088 6264 21140 6316
rect 23572 6400 23624 6452
rect 24032 6443 24084 6452
rect 24032 6409 24041 6443
rect 24041 6409 24075 6443
rect 24075 6409 24084 6443
rect 24032 6400 24084 6409
rect 25044 6443 25096 6452
rect 25044 6409 25053 6443
rect 25053 6409 25087 6443
rect 25087 6409 25096 6443
rect 25044 6400 25096 6409
rect 25136 6400 25188 6452
rect 27068 6443 27120 6452
rect 27068 6409 27077 6443
rect 27077 6409 27111 6443
rect 27111 6409 27120 6443
rect 27068 6400 27120 6409
rect 23940 6332 23992 6384
rect 21456 6196 21508 6248
rect 23756 6264 23808 6316
rect 27804 6332 27856 6384
rect 28540 6375 28592 6384
rect 28540 6341 28549 6375
rect 28549 6341 28583 6375
rect 28583 6341 28592 6375
rect 28540 6332 28592 6341
rect 37096 6332 37148 6384
rect 24768 6264 24820 6316
rect 19156 6128 19208 6180
rect 23112 6128 23164 6180
rect 24676 6196 24728 6248
rect 25320 6264 25372 6316
rect 26516 6264 26568 6316
rect 28816 6307 28868 6316
rect 28816 6273 28825 6307
rect 28825 6273 28859 6307
rect 28859 6273 28868 6307
rect 38016 6307 38068 6316
rect 28816 6264 28868 6273
rect 38016 6273 38025 6307
rect 38025 6273 38059 6307
rect 38059 6273 38068 6307
rect 38016 6264 38068 6273
rect 19892 6060 19944 6112
rect 23480 6060 23532 6112
rect 23848 6103 23900 6112
rect 23848 6069 23857 6103
rect 23857 6069 23891 6103
rect 23891 6069 23900 6103
rect 23848 6060 23900 6069
rect 36728 6103 36780 6112
rect 36728 6069 36737 6103
rect 36737 6069 36771 6103
rect 36771 6069 36780 6103
rect 36728 6060 36780 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 20260 5856 20312 5908
rect 22008 5856 22060 5908
rect 27804 5856 27856 5908
rect 2044 5652 2096 5704
rect 2780 5652 2832 5704
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4988 5652 5040 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 17408 5652 17460 5704
rect 18052 5720 18104 5772
rect 19340 5720 19392 5772
rect 20628 5763 20680 5772
rect 20628 5729 20637 5763
rect 20637 5729 20671 5763
rect 20671 5729 20680 5763
rect 20628 5720 20680 5729
rect 23572 5720 23624 5772
rect 17960 5652 18012 5704
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 18972 5652 19024 5704
rect 19432 5652 19484 5704
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 23848 5652 23900 5704
rect 37096 5763 37148 5772
rect 37096 5729 37105 5763
rect 37105 5729 37139 5763
rect 37139 5729 37148 5763
rect 37096 5720 37148 5729
rect 25228 5695 25280 5704
rect 25228 5661 25237 5695
rect 25237 5661 25271 5695
rect 25271 5661 25280 5695
rect 25228 5652 25280 5661
rect 25780 5652 25832 5704
rect 30380 5652 30432 5704
rect 34520 5652 34572 5704
rect 38108 5695 38160 5704
rect 38108 5661 38117 5695
rect 38117 5661 38151 5695
rect 38151 5661 38160 5695
rect 38108 5652 38160 5661
rect 3424 5584 3476 5636
rect 3056 5516 3108 5568
rect 16580 5516 16632 5568
rect 17132 5516 17184 5568
rect 19248 5516 19300 5568
rect 20076 5584 20128 5636
rect 37924 5627 37976 5636
rect 37924 5593 37933 5627
rect 37933 5593 37967 5627
rect 37967 5593 37976 5627
rect 37924 5584 37976 5593
rect 20812 5516 20864 5568
rect 23112 5516 23164 5568
rect 25872 5516 25924 5568
rect 25964 5559 26016 5568
rect 25964 5525 25973 5559
rect 25973 5525 26007 5559
rect 26007 5525 26016 5559
rect 25964 5516 26016 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 16028 5312 16080 5364
rect 18512 5312 18564 5364
rect 18604 5355 18656 5364
rect 18604 5321 18613 5355
rect 18613 5321 18647 5355
rect 18647 5321 18656 5355
rect 18604 5312 18656 5321
rect 20352 5312 20404 5364
rect 23940 5355 23992 5364
rect 23940 5321 23967 5355
rect 23967 5321 23992 5355
rect 23940 5312 23992 5321
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 36452 5312 36504 5364
rect 37924 5312 37976 5364
rect 3424 5287 3476 5296
rect 3424 5253 3433 5287
rect 3433 5253 3467 5287
rect 3467 5253 3476 5287
rect 3424 5244 3476 5253
rect 17132 5287 17184 5296
rect 17132 5253 17141 5287
rect 17141 5253 17175 5287
rect 17175 5253 17184 5287
rect 17132 5244 17184 5253
rect 17868 5244 17920 5296
rect 19340 5244 19392 5296
rect 23112 5244 23164 5296
rect 23572 5244 23624 5296
rect 25688 5244 25740 5296
rect 25872 5244 25924 5296
rect 3792 5176 3844 5228
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 16120 5219 16172 5228
rect 16120 5185 16129 5219
rect 16129 5185 16163 5219
rect 16163 5185 16172 5219
rect 16120 5176 16172 5185
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 15936 5108 15988 5160
rect 4068 5015 4120 5024
rect 4068 4981 4077 5015
rect 4077 4981 4111 5015
rect 4111 4981 4120 5015
rect 4068 4972 4120 4981
rect 5172 4972 5224 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 19984 5108 20036 5160
rect 20352 5040 20404 5092
rect 36636 5176 36688 5228
rect 23204 5151 23256 5160
rect 23204 5117 23213 5151
rect 23213 5117 23247 5151
rect 23247 5117 23256 5151
rect 23204 5108 23256 5117
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 28264 5108 28316 5160
rect 19432 4972 19484 5024
rect 22192 4972 22244 5024
rect 22376 4972 22428 5024
rect 23664 4972 23716 5024
rect 32588 4972 32640 5024
rect 34796 4972 34848 5024
rect 36636 4972 36688 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 16764 4768 16816 4820
rect 16856 4768 16908 4820
rect 17868 4811 17920 4820
rect 17868 4777 17877 4811
rect 17877 4777 17911 4811
rect 17911 4777 17920 4811
rect 17868 4768 17920 4777
rect 3056 4675 3108 4684
rect 3056 4641 3065 4675
rect 3065 4641 3099 4675
rect 3099 4641 3108 4675
rect 3056 4632 3108 4641
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 664 4496 716 4548
rect 2780 4496 2832 4548
rect 10784 4632 10836 4684
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 8944 4564 8996 4616
rect 9036 4564 9088 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 4160 4428 4212 4480
rect 11428 4428 11480 4480
rect 15936 4632 15988 4684
rect 16120 4632 16172 4684
rect 20352 4768 20404 4820
rect 22100 4768 22152 4820
rect 23204 4768 23256 4820
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 16580 4496 16632 4548
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 23296 4700 23348 4752
rect 21732 4632 21784 4684
rect 24768 4632 24820 4684
rect 26424 4632 26476 4684
rect 33140 4675 33192 4684
rect 33140 4641 33149 4675
rect 33149 4641 33183 4675
rect 33183 4641 33192 4675
rect 33140 4632 33192 4641
rect 37280 4632 37332 4684
rect 23388 4564 23440 4616
rect 19984 4496 20036 4548
rect 22100 4539 22152 4548
rect 22100 4505 22109 4539
rect 22109 4505 22143 4539
rect 22143 4505 22152 4539
rect 22100 4496 22152 4505
rect 23112 4496 23164 4548
rect 24492 4471 24544 4480
rect 24492 4437 24501 4471
rect 24501 4437 24535 4471
rect 24535 4437 24544 4471
rect 24492 4428 24544 4437
rect 31760 4564 31812 4616
rect 34704 4564 34756 4616
rect 25964 4496 26016 4548
rect 26240 4496 26292 4548
rect 32404 4539 32456 4548
rect 32404 4505 32413 4539
rect 32413 4505 32447 4539
rect 32447 4505 32456 4539
rect 32404 4496 32456 4505
rect 37556 4539 37608 4548
rect 37556 4505 37565 4539
rect 37565 4505 37599 4539
rect 37599 4505 37608 4539
rect 37556 4496 37608 4505
rect 25780 4428 25832 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 19984 4224 20036 4276
rect 22100 4224 22152 4276
rect 3424 4156 3476 4208
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 8300 4020 8352 4072
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 10876 4088 10928 4140
rect 18696 4088 18748 4140
rect 24492 4156 24544 4208
rect 20720 4131 20772 4140
rect 20720 4097 20729 4131
rect 20729 4097 20763 4131
rect 20763 4097 20772 4131
rect 20720 4088 20772 4097
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 22192 4020 22244 4072
rect 23204 4088 23256 4140
rect 24768 4131 24820 4140
rect 24768 4097 24777 4131
rect 24777 4097 24811 4131
rect 24811 4097 24820 4131
rect 25688 4131 25740 4140
rect 24768 4088 24820 4097
rect 25688 4097 25697 4131
rect 25697 4097 25731 4131
rect 25731 4097 25740 4131
rect 25688 4088 25740 4097
rect 25780 4131 25832 4140
rect 25780 4097 25789 4131
rect 25789 4097 25823 4131
rect 25823 4097 25832 4131
rect 25780 4088 25832 4097
rect 32588 4131 32640 4140
rect 23020 4063 23072 4072
rect 23020 4029 23029 4063
rect 23029 4029 23063 4063
rect 23063 4029 23072 4063
rect 23020 4020 23072 4029
rect 23480 4020 23532 4072
rect 6552 3952 6604 4004
rect 20076 3952 20128 4004
rect 21640 3952 21692 4004
rect 5908 3884 5960 3936
rect 6276 3884 6328 3936
rect 9220 3884 9272 3936
rect 10600 3884 10652 3936
rect 11244 3884 11296 3936
rect 13820 3884 13872 3936
rect 22376 3884 22428 3936
rect 32588 4097 32597 4131
rect 32597 4097 32631 4131
rect 32631 4097 32640 4131
rect 32588 4088 32640 4097
rect 36728 4131 36780 4140
rect 36728 4097 36737 4131
rect 36737 4097 36771 4131
rect 36771 4097 36780 4131
rect 37280 4131 37332 4140
rect 36728 4088 36780 4097
rect 37280 4097 37289 4131
rect 37289 4097 37323 4131
rect 37323 4097 37332 4131
rect 37280 4088 37332 4097
rect 38108 4131 38160 4140
rect 38108 4097 38117 4131
rect 38117 4097 38151 4131
rect 38151 4097 38160 4131
rect 38108 4088 38160 4097
rect 33416 4020 33468 4072
rect 33508 4063 33560 4072
rect 33508 4029 33517 4063
rect 33517 4029 33551 4063
rect 33551 4029 33560 4063
rect 35808 4063 35860 4072
rect 33508 4020 33560 4029
rect 35808 4029 35817 4063
rect 35817 4029 35851 4063
rect 35851 4029 35860 4063
rect 35808 4020 35860 4029
rect 37832 4020 37884 4072
rect 31208 3884 31260 3936
rect 33600 3884 33652 3936
rect 37924 3884 37976 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 8392 3680 8444 3732
rect 13360 3680 13412 3732
rect 23112 3723 23164 3732
rect 23112 3689 23121 3723
rect 23121 3689 23155 3723
rect 23155 3689 23164 3723
rect 23112 3680 23164 3689
rect 33416 3723 33468 3732
rect 33416 3689 33425 3723
rect 33425 3689 33459 3723
rect 33459 3689 33468 3723
rect 33416 3680 33468 3689
rect 37832 3723 37884 3732
rect 37832 3689 37841 3723
rect 37841 3689 37875 3723
rect 37875 3689 37884 3723
rect 37832 3680 37884 3689
rect 3424 3612 3476 3664
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6092 3544 6144 3596
rect 10968 3612 11020 3664
rect 1768 3476 1820 3528
rect 2964 3476 3016 3528
rect 6000 3476 6052 3528
rect 4160 3408 4212 3460
rect 4344 3408 4396 3460
rect 1952 3340 2004 3392
rect 3056 3340 3108 3392
rect 5080 3340 5132 3392
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 10784 3587 10836 3596
rect 10784 3553 10793 3587
rect 10793 3553 10827 3587
rect 10827 3553 10836 3587
rect 10784 3544 10836 3553
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 11428 3587 11480 3596
rect 11428 3553 11437 3587
rect 11437 3553 11471 3587
rect 11471 3553 11480 3587
rect 11428 3544 11480 3553
rect 14280 3544 14332 3596
rect 14556 3476 14608 3528
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 18972 3476 19024 3528
rect 32496 3612 32548 3664
rect 21180 3587 21232 3596
rect 21180 3553 21189 3587
rect 21189 3553 21223 3587
rect 21223 3553 21232 3587
rect 21180 3544 21232 3553
rect 22376 3587 22428 3596
rect 22376 3553 22385 3587
rect 22385 3553 22419 3587
rect 22419 3553 22428 3587
rect 22376 3544 22428 3553
rect 31208 3587 31260 3596
rect 31208 3553 31217 3587
rect 31217 3553 31251 3587
rect 31251 3553 31260 3587
rect 31208 3544 31260 3553
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 37924 3612 37976 3664
rect 36820 3587 36872 3596
rect 36820 3553 36829 3587
rect 36829 3553 36863 3587
rect 36863 3553 36872 3587
rect 36820 3544 36872 3553
rect 22560 3519 22612 3528
rect 22560 3485 22569 3519
rect 22569 3485 22603 3519
rect 22603 3485 22612 3519
rect 22560 3476 22612 3485
rect 23388 3476 23440 3528
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 24308 3408 24360 3460
rect 9128 3340 9180 3392
rect 14464 3340 14516 3392
rect 16856 3340 16908 3392
rect 19156 3340 19208 3392
rect 19432 3340 19484 3392
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 30748 3408 30800 3460
rect 33600 3476 33652 3528
rect 34704 3476 34756 3528
rect 37740 3519 37792 3528
rect 34428 3408 34480 3460
rect 37740 3485 37749 3519
rect 37749 3485 37783 3519
rect 37783 3485 37792 3519
rect 37740 3476 37792 3485
rect 37372 3408 37424 3460
rect 38200 3408 38252 3460
rect 35072 3340 35124 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4344 3179 4396 3188
rect 4344 3145 4353 3179
rect 4353 3145 4387 3179
rect 4387 3145 4396 3179
rect 4344 3136 4396 3145
rect 5632 3136 5684 3188
rect 16304 3136 16356 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 9220 3111 9272 3120
rect 9220 3077 9229 3111
rect 9229 3077 9263 3111
rect 9263 3077 9272 3111
rect 9220 3068 9272 3077
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 16856 3111 16908 3120
rect 16856 3077 16865 3111
rect 16865 3077 16899 3111
rect 16899 3077 16908 3111
rect 16856 3068 16908 3077
rect 19156 3111 19208 3120
rect 19156 3077 19165 3111
rect 19165 3077 19199 3111
rect 19199 3077 19208 3111
rect 19156 3068 19208 3077
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 4160 3000 4212 3052
rect 5080 3043 5132 3052
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 14280 3043 14332 3052
rect 13820 3000 13872 3009
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 4620 2932 4672 2984
rect 3884 2864 3936 2916
rect 6644 2932 6696 2984
rect 9680 2975 9732 2984
rect 9680 2941 9689 2975
rect 9689 2941 9723 2975
rect 9723 2941 9732 2975
rect 9680 2932 9732 2941
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 16672 2975 16724 2984
rect 16672 2941 16681 2975
rect 16681 2941 16715 2975
rect 16715 2941 16724 2975
rect 16672 2932 16724 2941
rect 18052 2932 18104 2984
rect 5448 2796 5500 2848
rect 6828 2796 6880 2848
rect 13544 2864 13596 2916
rect 16764 2864 16816 2916
rect 24308 3068 24360 3120
rect 22008 2975 22060 2984
rect 22008 2941 22017 2975
rect 22017 2941 22051 2975
rect 22051 2941 22060 2975
rect 22008 2932 22060 2941
rect 22468 2864 22520 2916
rect 21916 2796 21968 2848
rect 32404 3136 32456 3188
rect 32496 3136 32548 3188
rect 24768 3111 24820 3120
rect 24768 3077 24777 3111
rect 24777 3077 24811 3111
rect 24811 3077 24820 3111
rect 24768 3068 24820 3077
rect 35072 3111 35124 3120
rect 35072 3077 35081 3111
rect 35081 3077 35115 3111
rect 35115 3077 35124 3111
rect 35072 3068 35124 3077
rect 30748 3043 30800 3052
rect 30748 3009 30757 3043
rect 30757 3009 30791 3043
rect 30791 3009 30800 3043
rect 30748 3000 30800 3009
rect 31392 3043 31444 3052
rect 31392 3009 31401 3043
rect 31401 3009 31435 3043
rect 31435 3009 31444 3043
rect 31392 3000 31444 3009
rect 34796 3000 34848 3052
rect 37464 3000 37516 3052
rect 24584 2975 24636 2984
rect 24584 2941 24593 2975
rect 24593 2941 24627 2975
rect 24627 2941 24636 2975
rect 24584 2932 24636 2941
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 32128 2975 32180 2984
rect 32128 2941 32137 2975
rect 32137 2941 32171 2975
rect 32171 2941 32180 2975
rect 32128 2932 32180 2941
rect 35440 2975 35492 2984
rect 35440 2941 35449 2975
rect 35449 2941 35483 2975
rect 35483 2941 35492 2975
rect 35440 2932 35492 2941
rect 32220 2864 32272 2916
rect 34428 2796 34480 2848
rect 36544 2796 36596 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 13636 2592 13688 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 22008 2592 22060 2644
rect 22468 2635 22520 2644
rect 22468 2601 22477 2635
rect 22477 2601 22511 2635
rect 22511 2601 22520 2635
rect 22468 2592 22520 2601
rect 22560 2592 22612 2644
rect 24584 2592 24636 2644
rect 32128 2592 32180 2644
rect 37924 2635 37976 2644
rect 19432 2524 19484 2576
rect 31760 2524 31812 2576
rect 3056 2499 3108 2508
rect 3056 2465 3065 2499
rect 3065 2465 3099 2499
rect 3099 2465 3108 2499
rect 3056 2456 3108 2465
rect 4068 2456 4120 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 6000 2456 6052 2508
rect 6276 2456 6328 2508
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 6828 2499 6880 2508
rect 6828 2465 6837 2499
rect 6837 2465 6871 2499
rect 6871 2465 6880 2499
rect 6828 2456 6880 2465
rect 8392 2456 8444 2508
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 37924 2601 37933 2635
rect 37933 2601 37967 2635
rect 37967 2601 37976 2635
rect 37924 2592 37976 2601
rect 38016 2524 38068 2576
rect 36544 2499 36596 2508
rect 36544 2465 36553 2499
rect 36553 2465 36587 2499
rect 36587 2465 36596 2499
rect 36544 2456 36596 2465
rect 36728 2499 36780 2508
rect 36728 2465 36737 2499
rect 36737 2465 36771 2499
rect 36771 2465 36780 2499
rect 36728 2456 36780 2465
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 1400 2363 1452 2372
rect 1400 2329 1409 2363
rect 1409 2329 1443 2363
rect 1443 2329 1452 2363
rect 1400 2320 1452 2329
rect 9128 2363 9180 2372
rect 9128 2329 9137 2363
rect 9137 2329 9171 2363
rect 9171 2329 9180 2363
rect 9128 2320 9180 2329
rect 21548 2320 21600 2372
rect 34520 2388 34572 2440
rect 36912 2388 36964 2440
rect 35164 2320 35216 2372
rect 3240 2252 3292 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect -10 39200 102 40000
rect 634 39200 746 40000
rect 1278 39200 1390 40000
rect 1922 39200 2034 40000
rect 2566 39200 2678 40000
rect 3854 39200 3966 40000
rect 4498 39200 4610 40000
rect 5142 39200 5254 40000
rect 5786 39200 5898 40000
rect 6430 39200 6542 40000
rect 7074 39200 7186 40000
rect 7718 39200 7830 40000
rect 9006 39200 9118 40000
rect 9650 39200 9762 40000
rect 10294 39200 10406 40000
rect 10938 39200 11050 40000
rect 11582 39200 11694 40000
rect 12226 39200 12338 40000
rect 12870 39200 12982 40000
rect 14158 39200 14270 40000
rect 14802 39200 14914 40000
rect 15446 39200 15558 40000
rect 16090 39200 16202 40000
rect 16734 39200 16846 40000
rect 17378 39200 17490 40000
rect 18022 39200 18134 40000
rect 19310 39200 19422 40000
rect 19954 39200 20066 40000
rect 20598 39200 20710 40000
rect 21242 39200 21354 40000
rect 21886 39200 21998 40000
rect 22530 39200 22642 40000
rect 23174 39200 23286 40000
rect 24462 39200 24574 40000
rect 25106 39200 25218 40000
rect 25750 39200 25862 40000
rect 26394 39200 26506 40000
rect 27038 39200 27150 40000
rect 27682 39200 27794 40000
rect 28326 39200 28438 40000
rect 29614 39200 29726 40000
rect 30258 39200 30370 40000
rect 30902 39200 31014 40000
rect 31546 39200 31658 40000
rect 32190 39200 32302 40000
rect 32834 39200 32946 40000
rect 33478 39200 33590 40000
rect 34766 39200 34878 40000
rect 35410 39200 35522 40000
rect 36054 39200 36166 40000
rect 36698 39200 36810 40000
rect 37342 39200 37454 40000
rect 37986 39200 38098 40000
rect 38630 39200 38742 40000
rect 39274 39200 39386 40000
rect 1320 36242 1348 39200
rect 1582 37496 1638 37505
rect 1582 37431 1638 37440
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1412 36825 1440 37198
rect 1596 36854 1624 37431
rect 1964 37194 1992 39200
rect 2870 38856 2926 38865
rect 2870 38791 2926 38800
rect 2136 37256 2188 37262
rect 2136 37198 2188 37204
rect 1952 37188 2004 37194
rect 1952 37130 2004 37136
rect 2044 37120 2096 37126
rect 2044 37062 2096 37068
rect 2056 36922 2084 37062
rect 2044 36916 2096 36922
rect 2044 36858 2096 36864
rect 1584 36848 1636 36854
rect 1398 36816 1454 36825
rect 1584 36790 1636 36796
rect 1398 36751 1454 36760
rect 2148 36310 2176 37198
rect 2228 37120 2280 37126
rect 2228 37062 2280 37068
rect 2240 36854 2268 37062
rect 2228 36848 2280 36854
rect 2228 36790 2280 36796
rect 2136 36304 2188 36310
rect 2136 36246 2188 36252
rect 1308 36236 1360 36242
rect 1308 36178 1360 36184
rect 1768 35624 1820 35630
rect 1768 35566 1820 35572
rect 1780 34610 1808 35566
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1398 32056 1454 32065
rect 1398 31991 1454 32000
rect 1412 31890 1440 31991
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1872 25906 1900 26318
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 2148 21434 2176 36246
rect 2778 36136 2834 36145
rect 2778 36071 2834 36080
rect 2792 35630 2820 36071
rect 2228 35624 2280 35630
rect 2228 35566 2280 35572
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2240 34746 2268 35566
rect 2884 35154 2912 38791
rect 3056 37120 3108 37126
rect 3056 37062 3108 37068
rect 3068 36242 3096 37062
rect 3896 36854 3924 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 3884 36848 3936 36854
rect 3884 36790 3936 36796
rect 3424 36712 3476 36718
rect 3424 36654 3476 36660
rect 3056 36236 3108 36242
rect 3056 36178 3108 36184
rect 2964 36100 3016 36106
rect 2964 36042 3016 36048
rect 2872 35148 2924 35154
rect 2872 35090 2924 35096
rect 2872 35012 2924 35018
rect 2872 34954 2924 34960
rect 2884 34746 2912 34954
rect 2228 34740 2280 34746
rect 2228 34682 2280 34688
rect 2872 34740 2924 34746
rect 2872 34682 2924 34688
rect 2318 34640 2374 34649
rect 2318 34575 2320 34584
rect 2372 34575 2374 34584
rect 2320 34546 2372 34552
rect 2976 33522 3004 36042
rect 3240 35080 3292 35086
rect 3240 35022 3292 35028
rect 3252 34202 3280 35022
rect 3240 34196 3292 34202
rect 3240 34138 3292 34144
rect 3436 34134 3464 36654
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4632 36242 4660 37726
rect 9048 37618 9076 39200
rect 9048 37590 9168 37618
rect 5632 37256 5684 37262
rect 5632 37198 5684 37204
rect 6644 37256 6696 37262
rect 6644 37198 6696 37204
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 5540 36712 5592 36718
rect 5540 36654 5592 36660
rect 4620 36236 4672 36242
rect 4620 36178 4672 36184
rect 4620 36100 4672 36106
rect 4620 36042 4672 36048
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4632 35290 4660 36042
rect 5552 35834 5580 36654
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 4620 35284 4672 35290
rect 4620 35226 4672 35232
rect 5448 35012 5500 35018
rect 5448 34954 5500 34960
rect 3974 34776 4030 34785
rect 3974 34711 4030 34720
rect 3988 34542 4016 34711
rect 4712 34672 4764 34678
rect 4712 34614 4764 34620
rect 3608 34536 3660 34542
rect 3608 34478 3660 34484
rect 3792 34536 3844 34542
rect 3792 34478 3844 34484
rect 3976 34536 4028 34542
rect 3976 34478 4028 34484
rect 3424 34128 3476 34134
rect 3424 34070 3476 34076
rect 3620 33522 3648 34478
rect 3804 34202 3832 34478
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 3792 34196 3844 34202
rect 3792 34138 3844 34144
rect 2964 33516 3016 33522
rect 2964 33458 3016 33464
rect 3608 33516 3660 33522
rect 3608 33458 3660 33464
rect 3422 33416 3478 33425
rect 3422 33351 3424 33360
rect 3476 33351 3478 33360
rect 3424 33322 3476 33328
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4724 32842 4752 34614
rect 5264 33924 5316 33930
rect 5264 33866 5316 33872
rect 5276 33810 5304 33866
rect 5276 33782 5396 33810
rect 5368 33658 5396 33782
rect 5356 33652 5408 33658
rect 5356 33594 5408 33600
rect 5368 33454 5396 33594
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 4712 32836 4764 32842
rect 4712 32778 4764 32784
rect 3240 32224 3292 32230
rect 3240 32166 3292 32172
rect 3252 31890 3280 32166
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 3240 31884 3292 31890
rect 3240 31826 3292 31832
rect 3056 31748 3108 31754
rect 3056 31690 3108 31696
rect 3068 31482 3096 31690
rect 3056 31476 3108 31482
rect 3056 31418 3108 31424
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 2332 25265 2360 31282
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4158 29064 4214 29073
rect 4080 29022 4158 29050
rect 2870 25936 2926 25945
rect 2870 25871 2926 25880
rect 2884 25838 2912 25871
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2792 25498 2820 25774
rect 2780 25492 2832 25498
rect 2780 25434 2832 25440
rect 2318 25256 2374 25265
rect 2318 25191 2374 25200
rect 2148 21406 2268 21434
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 19922 1440 20878
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 19922 1624 20198
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 19825 1900 19858
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1688 18970 1716 19246
rect 1872 18970 1900 19246
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17746 1716 18022
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1964 17338 1992 17546
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2056 17202 2084 20402
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2148 19145 2176 19246
rect 2134 19136 2190 19145
rect 2134 19071 2190 19080
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16574 2084 17138
rect 2056 16546 2176 16574
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1400 14408 1452 14414
rect 1398 14376 1400 14385
rect 1452 14376 1454 14385
rect 1398 14311 1454 14320
rect 1872 13938 1900 14758
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2056 13530 2084 13806
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12306 1440 13262
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12306 1624 12582
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1952 11688 2004 11694
rect 2044 11688 2096 11694
rect 1952 11630 2004 11636
rect 2042 11656 2044 11665
rect 2096 11656 2098 11665
rect 1596 10674 1624 11630
rect 1964 11354 1992 11630
rect 2042 11591 2098 11600
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 9042 1440 9318
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1872 8945 1900 8978
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8634 1992 8842
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 7410 1808 7822
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1964 7002 1992 7278
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6322 1716 6734
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6390 1900 6598
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 2056 5710 2084 11086
rect 2148 8498 2176 16546
rect 2240 11150 2268 21406
rect 2332 18766 2360 25191
rect 4080 22094 4108 29022
rect 4158 28999 4214 29008
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4356 22642 4384 23054
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3988 22066 4108 22094
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 15570 3280 15846
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 3068 15162 3096 15370
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2792 14550 2820 14962
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 3068 14482 3096 14758
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13705 2820 13806
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2778 12336 2834 12345
rect 2778 12271 2780 12280
rect 2832 12271 2834 12280
rect 2780 12242 2832 12248
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2148 8022 2176 8434
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2792 7342 2820 7511
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2780 6248 2832 6254
rect 2778 6216 2780 6225
rect 2832 6216 2834 6225
rect 2778 6151 2834 6160
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4865 1808 5102
rect 1766 4856 1822 4865
rect 1766 4791 1822 4800
rect 2792 4554 2820 5646
rect 664 4548 716 4554
rect 664 4490 716 4496
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 676 800 704 4490
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1780 3058 1808 3470
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3126 1992 3334
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1412 2145 1440 2314
rect 1398 2136 1454 2145
rect 1398 2071 1454 2080
rect 2608 800 2636 4014
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2792 2825 2820 2926
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 2884 1465 2912 8366
rect 2976 6798 3004 12786
rect 3988 8974 4016 22066
rect 4632 21690 4660 23054
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4632 20482 4660 21626
rect 4540 20466 4660 20482
rect 4528 20460 4660 20466
rect 4580 20454 4660 20460
rect 4528 20402 4580 20408
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4632 19378 4660 20454
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4080 12850 4108 13466
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4080 8430 4108 9318
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8566 4384 8774
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 3988 7954 4016 8191
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4724 6914 4752 32778
rect 5080 31136 5132 31142
rect 5080 31078 5132 31084
rect 5172 31136 5224 31142
rect 5172 31078 5224 31084
rect 5092 30666 5120 31078
rect 5080 30660 5132 30666
rect 5080 30602 5132 30608
rect 5184 30258 5212 31078
rect 5172 30252 5224 30258
rect 5172 30194 5224 30200
rect 4804 30048 4856 30054
rect 4804 29990 4856 29996
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4816 29646 4844 29990
rect 4908 29850 4936 29990
rect 4896 29844 4948 29850
rect 4896 29786 4948 29792
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5092 13326 5120 13738
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4632 6886 4752 6914
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 3534 3004 6734
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 4690 3096 5510
rect 3252 4690 3280 5646
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3436 5302 3464 5578
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3804 5234 3832 5646
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3424 4208 3476 4214
rect 3422 4176 3424 4185
rect 3476 4176 3478 4185
rect 3422 4111 3478 4120
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 2964 3528 3016 3534
rect 3436 3505 3464 3606
rect 2964 3470 3016 3476
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3068 2514 3096 3334
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3252 800 3280 2246
rect 3896 800 3924 2858
rect 4080 2514 4108 4966
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4078 4200 4422
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4172 3058 4200 3402
rect 4356 3194 4384 3402
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4632 2990 4660 6886
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 4690 5028 5646
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4724 1714 4752 3538
rect 5092 3398 5120 13262
rect 5368 5234 5396 33390
rect 5460 29073 5488 34954
rect 5644 34202 5672 37198
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 6460 37120 6512 37126
rect 6460 37062 6512 37068
rect 5724 36916 5776 36922
rect 5724 36858 5776 36864
rect 5736 35737 5764 36858
rect 5828 36106 5856 37062
rect 6472 36786 6500 37062
rect 6656 36922 6684 37198
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 6644 36916 6696 36922
rect 6644 36858 6696 36864
rect 7194 36816 7250 36825
rect 6460 36780 6512 36786
rect 7194 36751 7196 36760
rect 6460 36722 6512 36728
rect 7248 36751 7250 36760
rect 7196 36722 7248 36728
rect 6472 36174 6500 36722
rect 6460 36168 6512 36174
rect 6460 36110 6512 36116
rect 5816 36100 5868 36106
rect 5816 36042 5868 36048
rect 5722 35728 5778 35737
rect 6472 35698 6500 36110
rect 7300 35766 7328 37062
rect 7760 36854 7788 37198
rect 7748 36848 7800 36854
rect 7748 36790 7800 36796
rect 8392 36712 8444 36718
rect 8392 36654 8444 36660
rect 9036 36712 9088 36718
rect 9036 36654 9088 36660
rect 7288 35760 7340 35766
rect 7288 35702 7340 35708
rect 8404 35698 8432 36654
rect 9048 36378 9076 36654
rect 9036 36372 9088 36378
rect 9036 36314 9088 36320
rect 8852 36168 8904 36174
rect 8852 36110 8904 36116
rect 5722 35663 5778 35672
rect 6460 35692 6512 35698
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 5736 34134 5764 35663
rect 6460 35634 6512 35640
rect 8392 35692 8444 35698
rect 8392 35634 8444 35640
rect 6000 35624 6052 35630
rect 6000 35566 6052 35572
rect 5816 35080 5868 35086
rect 5816 35022 5868 35028
rect 5724 34128 5776 34134
rect 5724 34070 5776 34076
rect 5828 33998 5856 35022
rect 6012 34202 6040 35566
rect 6472 35086 6500 35634
rect 7196 35624 7248 35630
rect 7196 35566 7248 35572
rect 6460 35080 6512 35086
rect 6460 35022 6512 35028
rect 6184 35012 6236 35018
rect 6184 34954 6236 34960
rect 6000 34196 6052 34202
rect 6000 34138 6052 34144
rect 5816 33992 5868 33998
rect 5816 33934 5868 33940
rect 5828 33522 5856 33934
rect 6012 33930 6040 34138
rect 6000 33924 6052 33930
rect 6000 33866 6052 33872
rect 5816 33516 5868 33522
rect 5816 33458 5868 33464
rect 5828 32910 5856 33458
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5724 32224 5776 32230
rect 5724 32166 5776 32172
rect 5736 31754 5764 32166
rect 6012 31754 6040 33866
rect 6196 31754 6224 34954
rect 6736 33516 6788 33522
rect 6736 33458 6788 33464
rect 6748 32502 6776 33458
rect 7208 33017 7236 35566
rect 8484 35080 8536 35086
rect 8484 35022 8536 35028
rect 8496 34542 8524 35022
rect 8864 35018 8892 36110
rect 9140 35834 9168 37590
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 9680 36644 9732 36650
rect 9680 36586 9732 36592
rect 9692 35834 9720 36586
rect 9784 36242 9812 37198
rect 9864 36372 9916 36378
rect 9864 36314 9916 36320
rect 9772 36236 9824 36242
rect 9772 36178 9824 36184
rect 9876 36122 9904 36314
rect 10336 36242 10364 39200
rect 10876 37188 10928 37194
rect 10876 37130 10928 37136
rect 10888 36922 10916 37130
rect 10876 36916 10928 36922
rect 10876 36858 10928 36864
rect 10508 36848 10560 36854
rect 10508 36790 10560 36796
rect 10416 36780 10468 36786
rect 10416 36722 10468 36728
rect 10428 36378 10456 36722
rect 10416 36372 10468 36378
rect 10416 36314 10468 36320
rect 10324 36236 10376 36242
rect 10324 36178 10376 36184
rect 9784 36106 9904 36122
rect 9772 36100 9904 36106
rect 9824 36094 9904 36100
rect 9956 36100 10008 36106
rect 9772 36042 9824 36048
rect 9956 36042 10008 36048
rect 9864 36032 9916 36038
rect 9864 35974 9916 35980
rect 9128 35828 9180 35834
rect 9128 35770 9180 35776
rect 9680 35828 9732 35834
rect 9680 35770 9732 35776
rect 9876 35698 9904 35974
rect 9968 35834 9996 36042
rect 9956 35828 10008 35834
rect 9956 35770 10008 35776
rect 9864 35692 9916 35698
rect 9864 35634 9916 35640
rect 8852 35012 8904 35018
rect 8852 34954 8904 34960
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 8484 34536 8536 34542
rect 8484 34478 8536 34484
rect 7470 33960 7526 33969
rect 7526 33904 7604 33912
rect 7470 33895 7472 33904
rect 7524 33884 7604 33904
rect 7472 33866 7524 33872
rect 7194 33008 7250 33017
rect 7194 32943 7250 32952
rect 6736 32496 6788 32502
rect 6736 32438 6788 32444
rect 6552 32360 6604 32366
rect 6552 32302 6604 32308
rect 6564 31822 6592 32302
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 5724 31748 5776 31754
rect 6012 31726 6132 31754
rect 6196 31726 6316 31754
rect 5724 31690 5776 31696
rect 5908 31340 5960 31346
rect 5908 31282 5960 31288
rect 5920 30598 5948 31282
rect 5908 30592 5960 30598
rect 5908 30534 5960 30540
rect 5920 30190 5948 30534
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5446 29064 5502 29073
rect 5446 28999 5502 29008
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5920 22098 5948 22374
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5460 21146 5488 21354
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5920 21010 5948 22034
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 6012 20806 6040 20878
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 7954 5672 8298
rect 5828 7954 5856 8910
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4690 5212 4966
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5184 4049 5212 4082
rect 5170 4040 5226 4049
rect 5170 3975 5226 3984
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 3058 5120 3334
rect 5644 3194 5672 6666
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5644 3058 5672 3130
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5460 2514 5488 2790
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 4540 1686 4752 1714
rect 4540 800 4568 1686
rect 5828 800 5856 4626
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5920 3602 5948 3878
rect 6104 3602 6132 31726
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6196 29034 6224 29582
rect 6184 29028 6236 29034
rect 6184 28970 6236 28976
rect 6196 27538 6224 28970
rect 6184 27532 6236 27538
rect 6184 27474 6236 27480
rect 6196 26994 6224 27474
rect 6184 26988 6236 26994
rect 6184 26930 6236 26936
rect 6196 25362 6224 26930
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 6288 22094 6316 31726
rect 6564 30802 6592 31758
rect 6748 31142 6776 32438
rect 6828 32428 6880 32434
rect 6828 32370 6880 32376
rect 7012 32428 7064 32434
rect 7012 32370 7064 32376
rect 6840 31482 6868 32370
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 6736 31136 6788 31142
rect 6736 31078 6788 31084
rect 7024 30802 7052 32370
rect 6552 30796 6604 30802
rect 6552 30738 6604 30744
rect 7012 30796 7064 30802
rect 7012 30738 7064 30744
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 7104 30660 7156 30666
rect 7104 30602 7156 30608
rect 6932 30394 6960 30602
rect 6920 30388 6972 30394
rect 6920 30330 6972 30336
rect 7116 30190 7144 30602
rect 7104 30184 7156 30190
rect 7104 30126 7156 30132
rect 7012 30116 7064 30122
rect 7012 30058 7064 30064
rect 7024 29646 7052 30058
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6564 27402 6592 27814
rect 7024 27606 7052 29582
rect 7116 28558 7144 30126
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 7012 27600 7064 27606
rect 7012 27542 7064 27548
rect 6552 27396 6604 27402
rect 6552 27338 6604 27344
rect 7116 27334 7144 28494
rect 7104 27328 7156 27334
rect 7104 27270 7156 27276
rect 6736 26920 6788 26926
rect 6736 26862 6788 26868
rect 6748 26586 6776 26862
rect 6736 26580 6788 26586
rect 6736 26522 6788 26528
rect 6552 25832 6604 25838
rect 6552 25774 6604 25780
rect 6564 25294 6592 25774
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6564 23730 6592 24006
rect 6932 23866 6960 24550
rect 7024 24206 7052 24754
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6368 23520 6420 23526
rect 6368 23462 6420 23468
rect 6380 23118 6408 23462
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6656 22642 6684 23666
rect 6736 23588 6788 23594
rect 6736 23530 6788 23536
rect 6748 22658 6776 23530
rect 6932 23526 6960 23802
rect 7024 23798 7052 24142
rect 7116 24138 7144 24686
rect 7104 24132 7156 24138
rect 7104 24074 7156 24080
rect 7012 23792 7064 23798
rect 7012 23734 7064 23740
rect 7116 23662 7144 24074
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6748 22642 6868 22658
rect 6552 22636 6604 22642
rect 6552 22578 6604 22584
rect 6644 22636 6696 22642
rect 6748 22636 6880 22642
rect 6748 22630 6828 22636
rect 6644 22578 6696 22584
rect 6828 22578 6880 22584
rect 6196 22066 6316 22094
rect 6196 20534 6224 22066
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6380 21690 6408 21966
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6380 21554 6408 21626
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6564 21146 6592 22578
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6656 21078 6684 21422
rect 6748 21350 6776 21966
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6748 20942 6776 21286
rect 6460 20936 6512 20942
rect 6736 20936 6788 20942
rect 6460 20878 6512 20884
rect 6656 20884 6736 20890
rect 6656 20878 6788 20884
rect 6184 20528 6236 20534
rect 6184 20470 6236 20476
rect 6472 19990 6500 20878
rect 6656 20862 6776 20878
rect 6656 20602 6684 20862
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6656 20058 6684 20402
rect 6748 20398 6776 20742
rect 6840 20534 6868 22578
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 7024 22030 7052 22510
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 7116 20534 7144 22170
rect 7208 22137 7236 32943
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7288 31884 7340 31890
rect 7288 31826 7340 31832
rect 7300 31414 7328 31826
rect 7392 31822 7420 32710
rect 7380 31816 7432 31822
rect 7380 31758 7432 31764
rect 7380 31680 7432 31686
rect 7380 31622 7432 31628
rect 7288 31408 7340 31414
rect 7288 31350 7340 31356
rect 7288 31272 7340 31278
rect 7288 31214 7340 31220
rect 7300 30666 7328 31214
rect 7288 30660 7340 30666
rect 7288 30602 7340 30608
rect 7392 30598 7420 31622
rect 7472 31204 7524 31210
rect 7472 31146 7524 31152
rect 7484 30734 7512 31146
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 7392 30326 7420 30534
rect 7380 30320 7432 30326
rect 7380 30262 7432 30268
rect 7484 30258 7512 30670
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7484 29714 7512 30194
rect 7576 29730 7604 33884
rect 8392 33312 8444 33318
rect 8392 33254 8444 33260
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 7656 32020 7708 32026
rect 7656 31962 7708 31968
rect 7668 31822 7696 31962
rect 7656 31816 7708 31822
rect 7656 31758 7708 31764
rect 7760 31482 7788 32846
rect 7852 31958 7880 32846
rect 8404 32502 8432 33254
rect 8496 32978 8524 34478
rect 9876 34202 9904 34546
rect 9956 34468 10008 34474
rect 9956 34410 10008 34416
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 9968 33998 9996 34410
rect 10140 34400 10192 34406
rect 10140 34342 10192 34348
rect 10152 34202 10180 34342
rect 10140 34196 10192 34202
rect 10140 34138 10192 34144
rect 9956 33992 10008 33998
rect 9956 33934 10008 33940
rect 10140 33856 10192 33862
rect 10140 33798 10192 33804
rect 10152 33386 10180 33798
rect 10232 33516 10284 33522
rect 10232 33458 10284 33464
rect 10140 33380 10192 33386
rect 10140 33322 10192 33328
rect 9128 33312 9180 33318
rect 9128 33254 9180 33260
rect 8484 32972 8536 32978
rect 8484 32914 8536 32920
rect 8496 32570 8524 32914
rect 9140 32842 9168 33254
rect 9128 32836 9180 32842
rect 9128 32778 9180 32784
rect 9772 32768 9824 32774
rect 10048 32768 10100 32774
rect 9824 32728 9996 32756
rect 9772 32710 9824 32716
rect 8484 32564 8536 32570
rect 8484 32506 8536 32512
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 8392 32224 8444 32230
rect 8392 32166 8444 32172
rect 7840 31952 7892 31958
rect 7840 31894 7892 31900
rect 7852 31822 7880 31894
rect 7840 31816 7892 31822
rect 8300 31816 8352 31822
rect 7840 31758 7892 31764
rect 8220 31776 8300 31804
rect 7748 31476 7800 31482
rect 7748 31418 7800 31424
rect 7748 31340 7800 31346
rect 7852 31328 7880 31758
rect 8220 31346 8248 31776
rect 8300 31758 8352 31764
rect 7800 31300 7880 31328
rect 7932 31340 7984 31346
rect 7748 31282 7800 31288
rect 7932 31282 7984 31288
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 7760 30938 7788 31282
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 7852 30598 7880 30738
rect 7944 30666 7972 31282
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 7932 30660 7984 30666
rect 7932 30602 7984 30608
rect 7840 30592 7892 30598
rect 7840 30534 7892 30540
rect 7472 29708 7524 29714
rect 7576 29702 7696 29730
rect 7472 29650 7524 29656
rect 7380 29232 7432 29238
rect 7380 29174 7432 29180
rect 7392 28626 7420 29174
rect 7484 29170 7512 29650
rect 7564 29640 7616 29646
rect 7564 29582 7616 29588
rect 7472 29164 7524 29170
rect 7472 29106 7524 29112
rect 7484 28966 7512 29106
rect 7576 29102 7604 29582
rect 7668 29152 7696 29702
rect 7852 29306 7880 30534
rect 8036 30394 8064 30670
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 8024 30116 8076 30122
rect 8024 30058 8076 30064
rect 8036 29578 8064 30058
rect 8024 29572 8076 29578
rect 8024 29514 8076 29520
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 7668 29124 7972 29152
rect 7564 29096 7616 29102
rect 7564 29038 7616 29044
rect 7472 28960 7524 28966
rect 7472 28902 7524 28908
rect 7748 28960 7800 28966
rect 7748 28902 7800 28908
rect 7380 28620 7432 28626
rect 7380 28562 7432 28568
rect 7392 28150 7420 28562
rect 7760 28490 7788 28902
rect 7748 28484 7800 28490
rect 7748 28426 7800 28432
rect 7380 28144 7432 28150
rect 7380 28086 7432 28092
rect 7288 28076 7340 28082
rect 7288 28018 7340 28024
rect 7300 25906 7328 28018
rect 7392 27402 7420 28086
rect 7760 28082 7788 28426
rect 7748 28076 7800 28082
rect 7748 28018 7800 28024
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7852 27470 7880 27814
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7380 27396 7432 27402
rect 7380 27338 7432 27344
rect 7380 27056 7432 27062
rect 7380 26998 7432 27004
rect 7392 26042 7420 26998
rect 7380 26036 7432 26042
rect 7380 25978 7432 25984
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7564 25220 7616 25226
rect 7564 25162 7616 25168
rect 7576 24410 7604 25162
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7668 23866 7696 24142
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7748 23792 7800 23798
rect 7748 23734 7800 23740
rect 7760 23186 7788 23734
rect 7748 23180 7800 23186
rect 7748 23122 7800 23128
rect 7760 22642 7788 23122
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7852 22710 7880 23054
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7194 22128 7250 22137
rect 7194 22063 7250 22072
rect 7576 21690 7604 22442
rect 7852 22250 7880 22646
rect 7668 22222 7880 22250
rect 7668 22166 7696 22222
rect 7656 22160 7708 22166
rect 7656 22102 7708 22108
rect 7838 22128 7894 22137
rect 7838 22063 7894 22072
rect 7852 21978 7880 22063
rect 7668 21950 7880 21978
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 6748 19854 6776 20334
rect 7116 19922 7144 20470
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 7116 19514 7144 19858
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6472 18970 6500 19314
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 7484 18766 7512 20198
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7668 15026 7696 21950
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7760 21486 7788 21830
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 7852 21078 7880 21490
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7852 19174 7880 20402
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7944 8498 7972 29124
rect 8036 27402 8064 29514
rect 8312 28082 8340 31078
rect 8404 30258 8432 32166
rect 9876 31822 9904 32302
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9876 31482 9904 31758
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9496 31408 9548 31414
rect 9496 31350 9548 31356
rect 9508 30938 9536 31350
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9496 30932 9548 30938
rect 9496 30874 9548 30880
rect 9600 30870 9628 31078
rect 9588 30864 9640 30870
rect 9588 30806 9640 30812
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 8392 30252 8444 30258
rect 8392 30194 8444 30200
rect 9680 30252 9732 30258
rect 9680 30194 9732 30200
rect 9128 29708 9180 29714
rect 9128 29650 9180 29656
rect 8576 29572 8628 29578
rect 8576 29514 8628 29520
rect 8588 29306 8616 29514
rect 8576 29300 8628 29306
rect 8576 29242 8628 29248
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 8496 28218 8524 29106
rect 9140 29102 9168 29650
rect 9128 29096 9180 29102
rect 9128 29038 9180 29044
rect 9692 28490 9720 30194
rect 9784 30054 9812 30670
rect 9864 30660 9916 30666
rect 9864 30602 9916 30608
rect 9876 30258 9904 30602
rect 9864 30252 9916 30258
rect 9864 30194 9916 30200
rect 9772 30048 9824 30054
rect 9772 29990 9824 29996
rect 9968 28994 9996 32728
rect 10048 32710 10100 32716
rect 10060 32434 10088 32710
rect 10048 32428 10100 32434
rect 10048 32370 10100 32376
rect 10244 31822 10272 33458
rect 10324 33312 10376 33318
rect 10324 33254 10376 33260
rect 10336 33114 10364 33254
rect 10324 33108 10376 33114
rect 10324 33050 10376 33056
rect 10336 32416 10364 33050
rect 10428 32994 10456 36314
rect 10520 35698 10548 36790
rect 10980 36650 11008 39200
rect 11520 37392 11572 37398
rect 11520 37334 11572 37340
rect 11624 37346 11652 39200
rect 11532 36786 11560 37334
rect 11624 37330 11744 37346
rect 11624 37324 11756 37330
rect 11624 37318 11704 37324
rect 11704 37266 11756 37272
rect 12164 37188 12216 37194
rect 12164 37130 12216 37136
rect 12072 36848 12124 36854
rect 12072 36790 12124 36796
rect 11520 36780 11572 36786
rect 11520 36722 11572 36728
rect 12084 36718 12112 36790
rect 11704 36712 11756 36718
rect 11704 36654 11756 36660
rect 12072 36712 12124 36718
rect 12072 36654 12124 36660
rect 10968 36644 11020 36650
rect 10968 36586 11020 36592
rect 10692 36576 10744 36582
rect 10692 36518 10744 36524
rect 10704 36038 10732 36518
rect 10692 36032 10744 36038
rect 10692 35974 10744 35980
rect 10704 35850 10732 35974
rect 10704 35822 11008 35850
rect 11716 35834 11744 36654
rect 12176 36174 12204 37130
rect 12268 36854 12296 39200
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 14188 37120 14240 37126
rect 14188 37062 14240 37068
rect 12728 36922 12756 37062
rect 12624 36916 12676 36922
rect 12624 36858 12676 36864
rect 12716 36916 12768 36922
rect 12716 36858 12768 36864
rect 12256 36848 12308 36854
rect 12256 36790 12308 36796
rect 12636 36378 12664 36858
rect 12624 36372 12676 36378
rect 12624 36314 12676 36320
rect 12164 36168 12216 36174
rect 12164 36110 12216 36116
rect 13544 36168 13596 36174
rect 13544 36110 13596 36116
rect 12176 35894 12204 36110
rect 12532 36100 12584 36106
rect 12532 36042 12584 36048
rect 13360 36100 13412 36106
rect 13360 36042 13412 36048
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12084 35866 12204 35894
rect 10508 35692 10560 35698
rect 10508 35634 10560 35640
rect 10520 33130 10548 35634
rect 10692 35148 10744 35154
rect 10692 35090 10744 35096
rect 10704 34950 10732 35090
rect 10784 35012 10836 35018
rect 10784 34954 10836 34960
rect 10600 34944 10652 34950
rect 10600 34886 10652 34892
rect 10692 34944 10744 34950
rect 10692 34886 10744 34892
rect 10612 34678 10640 34886
rect 10600 34672 10652 34678
rect 10600 34614 10652 34620
rect 10704 33386 10732 34886
rect 10796 34746 10824 34954
rect 10784 34740 10836 34746
rect 10784 34682 10836 34688
rect 10876 33516 10928 33522
rect 10876 33458 10928 33464
rect 10692 33380 10744 33386
rect 10692 33322 10744 33328
rect 10784 33312 10836 33318
rect 10784 33254 10836 33260
rect 10520 33102 10732 33130
rect 10428 32966 10548 32994
rect 10416 32836 10468 32842
rect 10416 32778 10468 32784
rect 10428 32570 10456 32778
rect 10416 32564 10468 32570
rect 10416 32506 10468 32512
rect 10416 32428 10468 32434
rect 10336 32388 10416 32416
rect 10416 32370 10468 32376
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10232 31816 10284 31822
rect 10232 31758 10284 31764
rect 10428 31754 10456 32166
rect 10416 31748 10468 31754
rect 10416 31690 10468 31696
rect 10048 31340 10100 31346
rect 10048 31282 10100 31288
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10060 30190 10088 31282
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10048 30184 10100 30190
rect 10048 30126 10100 30132
rect 9876 28966 9996 28994
rect 9876 28694 9904 28966
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9968 28490 9996 28698
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9956 28484 10008 28490
rect 9956 28426 10008 28432
rect 8944 28416 8996 28422
rect 8944 28358 8996 28364
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8116 28076 8168 28082
rect 8300 28076 8352 28082
rect 8168 28036 8300 28064
rect 8116 28018 8168 28024
rect 8300 28018 8352 28024
rect 8312 27953 8340 28018
rect 8024 27396 8076 27402
rect 8024 27338 8076 27344
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 8220 26450 8248 26862
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 8956 26314 8984 28358
rect 9312 28076 9364 28082
rect 9312 28018 9364 28024
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9140 26382 9168 27814
rect 9324 27470 9352 28018
rect 9692 28014 9720 28426
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 9876 28082 9904 28154
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9680 28008 9732 28014
rect 9680 27950 9732 27956
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9600 27538 9628 27814
rect 9692 27538 9720 27950
rect 9968 27538 9996 28426
rect 9588 27532 9640 27538
rect 9588 27474 9640 27480
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9312 27464 9364 27470
rect 9312 27406 9364 27412
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 9324 26382 9352 27270
rect 9692 27130 9720 27474
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9864 27056 9916 27062
rect 10060 27010 10088 30126
rect 10152 29322 10180 31078
rect 10244 30938 10272 31282
rect 10428 31142 10456 31690
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10428 30598 10456 31078
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10244 29510 10272 30194
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 10152 29294 10272 29322
rect 10140 29232 10192 29238
rect 10140 29174 10192 29180
rect 10152 28218 10180 29174
rect 10244 28558 10272 29294
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10140 28212 10192 28218
rect 10140 28154 10192 28160
rect 10244 28082 10272 28358
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 9864 26998 9916 27004
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 9128 25900 9180 25906
rect 9128 25842 9180 25848
rect 9140 25294 9168 25842
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 8220 24614 8248 25094
rect 8300 24880 8352 24886
rect 8300 24822 8352 24828
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8220 24206 8248 24550
rect 8312 24342 8340 24822
rect 8300 24336 8352 24342
rect 8300 24278 8352 24284
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8220 23798 8248 24142
rect 8312 23866 8340 24278
rect 8496 24274 8524 25094
rect 9140 24954 9168 25230
rect 9128 24948 9180 24954
rect 9128 24890 9180 24896
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9140 24410 9168 24754
rect 9220 24676 9272 24682
rect 9220 24618 9272 24624
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 9232 24206 9260 24618
rect 9692 24206 9720 25638
rect 9784 25498 9812 26726
rect 9876 26042 9904 26998
rect 9968 26982 10088 27010
rect 9968 26926 9996 26982
rect 9956 26920 10008 26926
rect 9956 26862 10008 26868
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 10244 25906 10272 28018
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 10336 26586 10364 26862
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10140 25900 10192 25906
rect 10140 25842 10192 25848
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9864 25220 9916 25226
rect 9864 25162 9916 25168
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9784 24206 9812 24550
rect 9876 24410 9904 25162
rect 10152 25158 10180 25842
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 10152 24818 10180 25094
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8128 22030 8156 23462
rect 8312 22658 8340 23802
rect 8496 23662 8524 24006
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8312 22642 8524 22658
rect 8588 22642 8616 24006
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8864 23322 8892 23666
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 8852 23316 8904 23322
rect 8852 23258 8904 23264
rect 8760 23044 8812 23050
rect 8760 22986 8812 22992
rect 8772 22778 8800 22986
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8300 22636 8524 22642
rect 8352 22630 8524 22636
rect 8300 22578 8352 22584
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8312 22234 8340 22374
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8404 21622 8432 22510
rect 8496 22506 8524 22630
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8864 22438 8892 23258
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8760 21956 8812 21962
rect 8760 21898 8812 21904
rect 8024 21616 8076 21622
rect 8024 21558 8076 21564
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8036 21418 8064 21558
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 8404 21146 8432 21558
rect 8772 21350 8800 21898
rect 8956 21486 8984 23054
rect 9416 22778 9444 23462
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 8128 20398 8156 20878
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8312 20466 8340 20810
rect 8772 20534 8800 21286
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8128 19922 8156 20334
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8956 19854 8984 21422
rect 9508 20534 9536 24074
rect 10152 23730 10180 24754
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 9692 22778 9720 23666
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 10152 22642 10180 23666
rect 10428 23322 10456 23666
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10428 23118 10456 23258
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10428 22234 10456 22442
rect 10416 22228 10468 22234
rect 10416 22170 10468 22176
rect 10230 22128 10286 22137
rect 10230 22063 10286 22072
rect 10520 22094 10548 32966
rect 10600 30932 10652 30938
rect 10600 30874 10652 30880
rect 10612 30394 10640 30874
rect 10600 30388 10652 30394
rect 10600 30330 10652 30336
rect 10704 26466 10732 33102
rect 10796 30802 10824 33254
rect 10888 33046 10916 33458
rect 10876 33040 10928 33046
rect 10876 32982 10928 32988
rect 10888 32366 10916 32982
rect 10876 32360 10928 32366
rect 10876 32302 10928 32308
rect 10888 31414 10916 32302
rect 10876 31408 10928 31414
rect 10876 31350 10928 31356
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10888 26586 10916 27406
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 10704 26438 10916 26466
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10612 22234 10640 23462
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10796 22642 10824 22918
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10704 22234 10732 22374
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10520 22066 10640 22094
rect 10244 22030 10272 22063
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 10244 20466 10272 21966
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 9600 19854 9628 20402
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 8680 19446 8708 19790
rect 8956 19446 8984 19790
rect 9036 19780 9088 19786
rect 9036 19722 9088 19728
rect 8668 19440 8720 19446
rect 8668 19382 8720 19388
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18290 8340 18566
rect 8680 18358 8708 19382
rect 9048 19378 9076 19722
rect 9784 19514 9812 20198
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9876 18834 9904 19450
rect 10336 19310 10364 19654
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9600 18426 9628 18702
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8036 17202 8064 17478
rect 8680 17270 8708 18294
rect 9692 17746 9720 18702
rect 10244 17746 10272 19178
rect 10336 18834 10364 19246
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 9692 17338 9720 17682
rect 9956 17604 10008 17610
rect 9956 17546 10008 17552
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 8668 17264 8720 17270
rect 8668 17206 8720 17212
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8680 16658 8708 17206
rect 9784 17202 9812 17478
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9968 17134 9996 17546
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8680 16182 8708 16594
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9232 16250 9260 16458
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 9416 16114 9444 16934
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9968 15638 9996 17070
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 10428 13802 10456 21354
rect 10520 21146 10548 21490
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 18222 10548 18566
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10520 17338 10548 18158
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6012 2514 6040 3470
rect 6288 2514 6316 3878
rect 6380 3058 6408 4966
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 7484 4146 7512 4558
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6564 2514 6592 3946
rect 8312 3738 8340 4014
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8404 3534 8432 3674
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6276 2508 6328 2514
rect 6276 2450 6328 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6656 2122 6684 2926
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2514 6868 2790
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 6472 2094 6684 2122
rect 6472 800 6500 2094
rect 8404 800 8432 2450
rect 8956 2446 8984 4558
rect 9048 3058 9076 4558
rect 9968 4146 9996 8434
rect 10612 6914 10640 22066
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10704 20992 10732 22034
rect 10796 22030 10824 22578
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10796 21690 10824 21966
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10784 21004 10836 21010
rect 10704 20964 10784 20992
rect 10784 20946 10836 20952
rect 10796 20330 10824 20946
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10796 19514 10824 19654
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10784 18896 10836 18902
rect 10704 18844 10784 18850
rect 10704 18838 10836 18844
rect 10704 18822 10824 18838
rect 10704 18766 10732 18822
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10704 17678 10732 18702
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 18426 10824 18566
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10704 16794 10732 17614
rect 10796 17338 10824 18362
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 15502 10824 16390
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10888 12434 10916 26438
rect 10980 21418 11008 35822
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11520 35624 11572 35630
rect 11520 35566 11572 35572
rect 11980 35624 12032 35630
rect 11980 35566 12032 35572
rect 11244 35488 11296 35494
rect 11244 35430 11296 35436
rect 11256 35086 11284 35430
rect 11244 35080 11296 35086
rect 11164 35040 11244 35068
rect 11060 34536 11112 34542
rect 11060 34478 11112 34484
rect 11072 33590 11100 34478
rect 11164 34082 11192 35040
rect 11244 35022 11296 35028
rect 11164 34066 11284 34082
rect 11152 34060 11284 34066
rect 11204 34054 11284 34060
rect 11152 34002 11204 34008
rect 11152 33924 11204 33930
rect 11152 33866 11204 33872
rect 11060 33584 11112 33590
rect 11060 33526 11112 33532
rect 11164 33454 11192 33866
rect 11152 33448 11204 33454
rect 11152 33390 11204 33396
rect 11256 33114 11284 34054
rect 11532 33386 11560 35566
rect 11992 35290 12020 35566
rect 11980 35284 12032 35290
rect 11980 35226 12032 35232
rect 11980 35012 12032 35018
rect 11980 34954 12032 34960
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11888 34944 11940 34950
rect 11888 34886 11940 34892
rect 11716 34610 11744 34886
rect 11900 34678 11928 34886
rect 11888 34672 11940 34678
rect 11888 34614 11940 34620
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 11992 34406 12020 34954
rect 12084 34542 12112 35866
rect 12452 35086 12480 35974
rect 12544 35766 12572 36042
rect 12532 35760 12584 35766
rect 12532 35702 12584 35708
rect 12532 35284 12584 35290
rect 12532 35226 12584 35232
rect 12164 35080 12216 35086
rect 12164 35022 12216 35028
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 12176 34610 12204 35022
rect 12544 35018 12572 35226
rect 13372 35086 13400 36042
rect 13556 35494 13584 36110
rect 14200 36106 14228 37062
rect 16132 36786 16160 37266
rect 17684 37256 17736 37262
rect 17684 37198 17736 37204
rect 17696 36786 17724 37198
rect 16120 36780 16172 36786
rect 16120 36722 16172 36728
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 17040 36712 17092 36718
rect 17040 36654 17092 36660
rect 16948 36576 17000 36582
rect 16948 36518 17000 36524
rect 16304 36236 16356 36242
rect 16304 36178 16356 36184
rect 14188 36100 14240 36106
rect 14188 36042 14240 36048
rect 15568 36100 15620 36106
rect 15568 36042 15620 36048
rect 14096 36032 14148 36038
rect 14096 35974 14148 35980
rect 14108 35698 14136 35974
rect 15580 35834 15608 36042
rect 15660 36032 15712 36038
rect 15660 35974 15712 35980
rect 15568 35828 15620 35834
rect 15568 35770 15620 35776
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 14372 35692 14424 35698
rect 14372 35634 14424 35640
rect 14464 35692 14516 35698
rect 14464 35634 14516 35640
rect 15108 35692 15160 35698
rect 15108 35634 15160 35640
rect 15292 35692 15344 35698
rect 15292 35634 15344 35640
rect 13820 35624 13872 35630
rect 13820 35566 13872 35572
rect 13544 35488 13596 35494
rect 13544 35430 13596 35436
rect 13636 35488 13688 35494
rect 13636 35430 13688 35436
rect 13556 35086 13584 35430
rect 13360 35080 13412 35086
rect 13360 35022 13412 35028
rect 13544 35080 13596 35086
rect 13544 35022 13596 35028
rect 12532 35012 12584 35018
rect 12532 34954 12584 34960
rect 12716 35012 12768 35018
rect 12716 34954 12768 34960
rect 12164 34604 12216 34610
rect 12164 34546 12216 34552
rect 12072 34536 12124 34542
rect 12072 34478 12124 34484
rect 11980 34400 12032 34406
rect 11980 34342 12032 34348
rect 11796 34196 11848 34202
rect 11796 34138 11848 34144
rect 11808 34082 11836 34138
rect 11716 34054 11836 34082
rect 11716 33862 11744 34054
rect 11992 33998 12020 34342
rect 12544 33998 12572 34954
rect 12728 34746 12756 34954
rect 12716 34740 12768 34746
rect 12716 34682 12768 34688
rect 13556 34474 13584 35022
rect 13648 34950 13676 35430
rect 13832 34950 13860 35566
rect 14108 35154 14136 35634
rect 14384 35494 14412 35634
rect 14372 35488 14424 35494
rect 14372 35430 14424 35436
rect 14476 35222 14504 35634
rect 14464 35216 14516 35222
rect 14464 35158 14516 35164
rect 14096 35148 14148 35154
rect 14096 35090 14148 35096
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 13636 34944 13688 34950
rect 13636 34886 13688 34892
rect 13820 34944 13872 34950
rect 13820 34886 13872 34892
rect 13176 34468 13228 34474
rect 13176 34410 13228 34416
rect 13544 34468 13596 34474
rect 13544 34410 13596 34416
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 11704 33856 11756 33862
rect 11704 33798 11756 33804
rect 11808 33590 11836 33934
rect 12624 33924 12676 33930
rect 12624 33866 12676 33872
rect 11888 33856 11940 33862
rect 12636 33833 12664 33866
rect 13084 33856 13136 33862
rect 11888 33798 11940 33804
rect 12622 33824 12678 33833
rect 11796 33584 11848 33590
rect 11796 33526 11848 33532
rect 11520 33380 11572 33386
rect 11520 33322 11572 33328
rect 11244 33108 11296 33114
rect 11244 33050 11296 33056
rect 11532 32978 11560 33322
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11900 32910 11928 33798
rect 13084 33798 13136 33804
rect 12622 33759 12678 33768
rect 12808 33584 12860 33590
rect 12808 33526 12860 33532
rect 12348 33448 12400 33454
rect 12348 33390 12400 33396
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11888 32904 11940 32910
rect 11888 32846 11940 32852
rect 11060 32496 11112 32502
rect 11060 32438 11112 32444
rect 11072 32298 11100 32438
rect 11060 32292 11112 32298
rect 11060 32234 11112 32240
rect 11072 31958 11100 32234
rect 11624 32230 11652 32846
rect 11796 32768 11848 32774
rect 11796 32710 11848 32716
rect 11808 32434 11836 32710
rect 11704 32428 11756 32434
rect 11704 32370 11756 32376
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11612 32224 11664 32230
rect 11612 32166 11664 32172
rect 11060 31952 11112 31958
rect 11112 31900 11284 31906
rect 11060 31894 11284 31900
rect 11072 31878 11284 31894
rect 11060 31816 11112 31822
rect 11060 31758 11112 31764
rect 11072 31482 11100 31758
rect 11060 31476 11112 31482
rect 11060 31418 11112 31424
rect 11152 30184 11204 30190
rect 11152 30126 11204 30132
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 11072 29238 11100 29650
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 11164 28694 11192 30126
rect 11256 29170 11284 31878
rect 11624 31754 11652 32166
rect 11716 32026 11744 32370
rect 11808 32026 11836 32370
rect 11704 32020 11756 32026
rect 11704 31962 11756 31968
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11440 31726 11652 31754
rect 11440 30122 11468 31726
rect 11520 31408 11572 31414
rect 11520 31350 11572 31356
rect 11532 30258 11560 31350
rect 11612 31272 11664 31278
rect 11612 31214 11664 31220
rect 11624 30734 11652 31214
rect 11716 31142 11744 31826
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 11716 30870 11744 31078
rect 11704 30864 11756 30870
rect 11704 30806 11756 30812
rect 11612 30728 11664 30734
rect 11900 30682 11928 32846
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 12176 31822 12204 32302
rect 12164 31816 12216 31822
rect 12164 31758 12216 31764
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 11612 30670 11664 30676
rect 11808 30654 11928 30682
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11428 30116 11480 30122
rect 11428 30058 11480 30064
rect 11532 30054 11560 30194
rect 11808 30138 11836 30654
rect 11888 30592 11940 30598
rect 11886 30560 11888 30569
rect 11940 30560 11942 30569
rect 11886 30495 11942 30504
rect 11900 30258 11928 30495
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 11612 30116 11664 30122
rect 11808 30110 11928 30138
rect 11612 30058 11664 30064
rect 11520 30048 11572 30054
rect 11520 29990 11572 29996
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 11348 28762 11376 29582
rect 11428 29572 11480 29578
rect 11428 29514 11480 29520
rect 11336 28756 11388 28762
rect 11336 28698 11388 28704
rect 11440 28694 11468 29514
rect 11532 29306 11560 29990
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 11428 28688 11480 28694
rect 11428 28630 11480 28636
rect 11440 28014 11468 28630
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 11624 27130 11652 30058
rect 11796 30048 11848 30054
rect 11796 29990 11848 29996
rect 11808 29170 11836 29990
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11716 27674 11744 28018
rect 11704 27668 11756 27674
rect 11704 27610 11756 27616
rect 11900 27554 11928 30110
rect 11992 30054 12020 30670
rect 12072 30592 12124 30598
rect 12072 30534 12124 30540
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 12084 29578 12112 30534
rect 12176 30326 12204 31078
rect 12268 30598 12296 32370
rect 12360 31346 12388 33390
rect 12820 32570 12848 33526
rect 12900 33448 12952 33454
rect 12900 33390 12952 33396
rect 12912 33114 12940 33390
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 13096 32910 13124 33798
rect 13084 32904 13136 32910
rect 13084 32846 13136 32852
rect 12808 32564 12860 32570
rect 12808 32506 12860 32512
rect 13084 32564 13136 32570
rect 13084 32506 13136 32512
rect 12992 32496 13044 32502
rect 12992 32438 13044 32444
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 13004 31278 13032 32438
rect 12716 31272 12768 31278
rect 12716 31214 12768 31220
rect 12992 31272 13044 31278
rect 12992 31214 13044 31220
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12256 30592 12308 30598
rect 12256 30534 12308 30540
rect 12164 30320 12216 30326
rect 12164 30262 12216 30268
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 11980 29096 12032 29102
rect 11980 29038 12032 29044
rect 11992 28994 12020 29038
rect 12176 28994 12204 30262
rect 12360 30258 12388 31078
rect 12728 30802 12756 31214
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 13004 30734 13032 31214
rect 12808 30728 12860 30734
rect 12992 30728 13044 30734
rect 12808 30670 12860 30676
rect 12912 30688 12992 30716
rect 12820 30394 12848 30670
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 12256 30184 12308 30190
rect 12256 30126 12308 30132
rect 12268 29578 12296 30126
rect 12360 29782 12388 30194
rect 12532 30184 12584 30190
rect 12584 30144 12664 30172
rect 12532 30126 12584 30132
rect 12636 29782 12664 30144
rect 12912 29866 12940 30688
rect 12992 30670 13044 30676
rect 12820 29850 12940 29866
rect 12808 29844 12940 29850
rect 12860 29838 12940 29844
rect 12808 29786 12860 29792
rect 12348 29776 12400 29782
rect 12348 29718 12400 29724
rect 12624 29776 12676 29782
rect 12624 29718 12676 29724
rect 12636 29646 12664 29718
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 12268 29481 12296 29514
rect 12440 29504 12492 29510
rect 12254 29472 12310 29481
rect 12440 29446 12492 29452
rect 12254 29407 12310 29416
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12268 29170 12296 29242
rect 12452 29170 12480 29446
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 11992 28966 12204 28994
rect 11992 28490 12020 28966
rect 12636 28626 12664 29582
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12912 29306 12940 29446
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 13004 29170 13032 29582
rect 12992 29164 13044 29170
rect 12992 29106 13044 29112
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 11980 28484 12032 28490
rect 11980 28426 12032 28432
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 12636 28014 12664 28358
rect 12728 28082 12756 28358
rect 12808 28144 12860 28150
rect 12808 28086 12860 28092
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12440 27872 12492 27878
rect 12440 27814 12492 27820
rect 11808 27526 11928 27554
rect 12256 27600 12308 27606
rect 12452 27554 12480 27814
rect 12308 27548 12480 27554
rect 12256 27542 12480 27548
rect 12268 27526 12480 27542
rect 12728 27538 12756 28018
rect 12820 27674 12848 28086
rect 13096 28082 13124 32506
rect 13188 32026 13216 34410
rect 13832 34066 13860 34886
rect 13924 34678 13952 35022
rect 14108 34678 14136 35090
rect 14464 35012 14516 35018
rect 14464 34954 14516 34960
rect 14188 34740 14240 34746
rect 14188 34682 14240 34688
rect 13912 34672 13964 34678
rect 13912 34614 13964 34620
rect 14096 34672 14148 34678
rect 14096 34614 14148 34620
rect 13912 34400 13964 34406
rect 13964 34360 14136 34388
rect 13912 34342 13964 34348
rect 13820 34060 13872 34066
rect 13820 34002 13872 34008
rect 13268 33992 13320 33998
rect 13320 33952 13400 33980
rect 13268 33934 13320 33940
rect 13268 33856 13320 33862
rect 13268 33798 13320 33804
rect 13176 32020 13228 32026
rect 13176 31962 13228 31968
rect 13280 31754 13308 33798
rect 13372 33454 13400 33952
rect 13360 33448 13412 33454
rect 13360 33390 13412 33396
rect 13372 32230 13400 33390
rect 14004 32904 14056 32910
rect 14004 32846 14056 32852
rect 13360 32224 13412 32230
rect 13360 32166 13412 32172
rect 14016 31890 14044 32846
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13268 31748 13320 31754
rect 13268 31690 13320 31696
rect 13280 30326 13308 31690
rect 13360 31136 13412 31142
rect 13360 31078 13412 31084
rect 13372 30734 13400 31078
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13268 30320 13320 30326
rect 13268 30262 13320 30268
rect 13372 29696 13400 30670
rect 13452 30320 13504 30326
rect 13452 30262 13504 30268
rect 13464 29850 13492 30262
rect 13452 29844 13504 29850
rect 13452 29786 13504 29792
rect 13452 29708 13504 29714
rect 13372 29668 13452 29696
rect 13452 29650 13504 29656
rect 13556 28082 13584 31758
rect 14016 30258 14044 31826
rect 14108 30870 14136 34360
rect 14200 33930 14228 34682
rect 14280 34604 14332 34610
rect 14280 34546 14332 34552
rect 14188 33924 14240 33930
rect 14188 33866 14240 33872
rect 14292 33454 14320 34546
rect 14372 34400 14424 34406
rect 14372 34342 14424 34348
rect 14384 33930 14412 34342
rect 14476 34202 14504 34954
rect 15120 34746 15148 35634
rect 15304 35290 15332 35634
rect 15292 35284 15344 35290
rect 15292 35226 15344 35232
rect 15292 35080 15344 35086
rect 15292 35022 15344 35028
rect 15200 34944 15252 34950
rect 15200 34886 15252 34892
rect 15108 34740 15160 34746
rect 15108 34682 15160 34688
rect 15212 34474 15240 34886
rect 15304 34542 15332 35022
rect 15384 35012 15436 35018
rect 15384 34954 15436 34960
rect 15396 34610 15424 34954
rect 15476 34944 15528 34950
rect 15476 34886 15528 34892
rect 15384 34604 15436 34610
rect 15384 34546 15436 34552
rect 15488 34542 15516 34886
rect 15292 34536 15344 34542
rect 15292 34478 15344 34484
rect 15476 34536 15528 34542
rect 15476 34478 15528 34484
rect 15200 34468 15252 34474
rect 15200 34410 15252 34416
rect 15108 34400 15160 34406
rect 15108 34342 15160 34348
rect 14464 34196 14516 34202
rect 14464 34138 14516 34144
rect 15120 34066 15148 34342
rect 15108 34060 15160 34066
rect 15108 34002 15160 34008
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 15200 33856 15252 33862
rect 15200 33798 15252 33804
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14280 33448 14332 33454
rect 14280 33390 14332 33396
rect 14292 33046 14320 33390
rect 14280 33040 14332 33046
rect 14280 32982 14332 32988
rect 14188 32768 14240 32774
rect 14188 32710 14240 32716
rect 14096 30864 14148 30870
rect 14096 30806 14148 30812
rect 14200 30802 14228 32710
rect 14280 31408 14332 31414
rect 14280 31350 14332 31356
rect 14188 30796 14240 30802
rect 14188 30738 14240 30744
rect 14188 30388 14240 30394
rect 14188 30330 14240 30336
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13648 29782 13676 29990
rect 13636 29776 13688 29782
rect 13636 29718 13688 29724
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 13648 29481 13676 29582
rect 13634 29472 13690 29481
rect 13634 29407 13690 29416
rect 13648 28150 13676 29407
rect 13832 29170 13860 29990
rect 14200 29578 14228 30330
rect 14188 29572 14240 29578
rect 14188 29514 14240 29520
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 14292 28218 14320 31350
rect 14568 31210 14596 33594
rect 15212 33590 15240 33798
rect 15304 33590 15332 34478
rect 15384 34060 15436 34066
rect 15384 34002 15436 34008
rect 15200 33584 15252 33590
rect 15200 33526 15252 33532
rect 15292 33584 15344 33590
rect 15292 33526 15344 33532
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 14648 33108 14700 33114
rect 14648 33050 14700 33056
rect 14660 32842 14688 33050
rect 15304 32910 15332 33390
rect 15396 32978 15424 34002
rect 15384 32972 15436 32978
rect 15384 32914 15436 32920
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 14648 32836 14700 32842
rect 14648 32778 14700 32784
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 14372 31204 14424 31210
rect 14372 31146 14424 31152
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 14384 29238 14412 31146
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14372 28960 14424 28966
rect 14372 28902 14424 28908
rect 14384 28490 14412 28902
rect 14476 28626 14504 30670
rect 14660 29170 14688 32778
rect 15212 32570 15240 32778
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 15304 32502 15332 32846
rect 15396 32570 15424 32914
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15488 32502 15516 34478
rect 15568 34468 15620 34474
rect 15568 34410 15620 34416
rect 15580 33833 15608 34410
rect 15672 33930 15700 35974
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 15948 35154 15976 35634
rect 16316 35601 16344 36178
rect 16396 36168 16448 36174
rect 16396 36110 16448 36116
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16408 35698 16436 36110
rect 16396 35692 16448 35698
rect 16396 35634 16448 35640
rect 16302 35592 16358 35601
rect 16302 35527 16358 35536
rect 16212 35216 16264 35222
rect 16212 35158 16264 35164
rect 15936 35148 15988 35154
rect 15936 35090 15988 35096
rect 16224 34746 16252 35158
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 16316 34202 16344 35022
rect 16212 34196 16264 34202
rect 16212 34138 16264 34144
rect 16304 34196 16356 34202
rect 16304 34138 16356 34144
rect 16224 33946 16252 34138
rect 16408 34066 16436 35634
rect 16396 34060 16448 34066
rect 16396 34002 16448 34008
rect 15660 33924 15712 33930
rect 16224 33918 16436 33946
rect 15660 33866 15712 33872
rect 15566 33824 15622 33833
rect 15566 33759 15622 33768
rect 15292 32496 15344 32502
rect 15292 32438 15344 32444
rect 15476 32496 15528 32502
rect 15476 32438 15528 32444
rect 15304 32042 15332 32438
rect 15580 32434 15608 33759
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 15212 32014 15332 32042
rect 15212 31822 15240 32014
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15016 31816 15068 31822
rect 15016 31758 15068 31764
rect 15200 31816 15252 31822
rect 15200 31758 15252 31764
rect 15028 31346 15056 31758
rect 15016 31340 15068 31346
rect 15016 31282 15068 31288
rect 14740 30660 14792 30666
rect 14740 30602 14792 30608
rect 14752 30394 14780 30602
rect 15028 30598 15056 31282
rect 15016 30592 15068 30598
rect 15304 30546 15332 31894
rect 15016 30534 15068 30540
rect 14740 30388 14792 30394
rect 14740 30330 14792 30336
rect 14740 30252 14792 30258
rect 14740 30194 14792 30200
rect 14752 29646 14780 30194
rect 15028 29646 15056 30534
rect 15212 30518 15332 30546
rect 15212 30326 15240 30518
rect 15396 30326 15424 32370
rect 15476 31136 15528 31142
rect 15476 31078 15528 31084
rect 15200 30320 15252 30326
rect 15200 30262 15252 30268
rect 15384 30320 15436 30326
rect 15384 30262 15436 30268
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15304 30138 15332 30194
rect 15488 30190 15516 31078
rect 15476 30184 15528 30190
rect 15304 30110 15424 30138
rect 15476 30126 15528 30132
rect 15108 29708 15160 29714
rect 15108 29650 15160 29656
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14752 29238 14780 29582
rect 14740 29232 14792 29238
rect 14740 29174 14792 29180
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14924 29028 14976 29034
rect 14924 28970 14976 28976
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 14372 28484 14424 28490
rect 14372 28426 14424 28432
rect 14476 28218 14504 28562
rect 14280 28212 14332 28218
rect 14280 28154 14332 28160
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 12900 28076 12952 28082
rect 12900 28018 12952 28024
rect 13084 28076 13136 28082
rect 13084 28018 13136 28024
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 14832 28076 14884 28082
rect 14832 28018 14884 28024
rect 12912 27878 12940 28018
rect 14844 27878 14872 28018
rect 14936 27878 14964 28970
rect 15028 27962 15056 29582
rect 15120 29102 15148 29650
rect 15396 29578 15424 30110
rect 15384 29572 15436 29578
rect 15384 29514 15436 29520
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 15108 29096 15160 29102
rect 15108 29038 15160 29044
rect 15120 28150 15148 29038
rect 15304 28150 15332 29174
rect 15396 28626 15424 29514
rect 15580 29306 15608 32370
rect 15660 31816 15712 31822
rect 15660 31758 15712 31764
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 15672 31346 15700 31758
rect 16316 31634 16344 31758
rect 16224 31606 16344 31634
rect 16028 31476 16080 31482
rect 16028 31418 16080 31424
rect 15660 31340 15712 31346
rect 15660 31282 15712 31288
rect 15752 30864 15804 30870
rect 15752 30806 15804 30812
rect 15660 30184 15712 30190
rect 15660 30126 15712 30132
rect 15672 29646 15700 30126
rect 15764 29850 15792 30806
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15764 29306 15792 29786
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15568 29300 15620 29306
rect 15568 29242 15620 29248
rect 15752 29300 15804 29306
rect 15752 29242 15804 29248
rect 15844 29232 15896 29238
rect 15844 29174 15896 29180
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15108 28144 15160 28150
rect 15108 28086 15160 28092
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 15028 27934 15148 27962
rect 15120 27878 15148 27934
rect 12900 27872 12952 27878
rect 12900 27814 12952 27820
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 14832 27872 14884 27878
rect 14832 27814 14884 27820
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 15108 27872 15160 27878
rect 15108 27814 15160 27820
rect 13096 27674 13124 27814
rect 12808 27668 12860 27674
rect 12808 27610 12860 27616
rect 13084 27668 13136 27674
rect 13084 27610 13136 27616
rect 14464 27600 14516 27606
rect 14464 27542 14516 27548
rect 12716 27532 12768 27538
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11624 26874 11652 27066
rect 11624 26846 11744 26874
rect 11716 26790 11744 26846
rect 11612 26784 11664 26790
rect 11612 26726 11664 26732
rect 11704 26784 11756 26790
rect 11704 26726 11756 26732
rect 11624 25906 11652 26726
rect 11808 26058 11836 27526
rect 12716 27474 12768 27480
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 13544 27464 13596 27470
rect 13544 27406 13596 27412
rect 11900 27130 11928 27406
rect 11888 27124 11940 27130
rect 11888 27066 11940 27072
rect 11900 26994 11928 27066
rect 13556 27062 13584 27406
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 13544 27056 13596 27062
rect 13544 26998 13596 27004
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 14108 26926 14136 27270
rect 14476 27130 14504 27542
rect 14844 27538 14872 27814
rect 14936 27606 14964 27814
rect 14924 27600 14976 27606
rect 14924 27542 14976 27548
rect 14832 27532 14884 27538
rect 14832 27474 14884 27480
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14280 27056 14332 27062
rect 14280 26998 14332 27004
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 11808 26030 11928 26058
rect 11796 25968 11848 25974
rect 11796 25910 11848 25916
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11624 25362 11652 25842
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11072 24682 11100 25230
rect 11060 24676 11112 24682
rect 11060 24618 11112 24624
rect 11624 24206 11652 25298
rect 11808 24954 11836 25910
rect 11900 25294 11928 26030
rect 11992 25498 12020 26318
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 12084 25974 12112 26182
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11808 24834 11836 24890
rect 11716 24806 11836 24834
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11520 24132 11572 24138
rect 11520 24074 11572 24080
rect 11532 23866 11560 24074
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11624 23798 11652 24142
rect 11612 23792 11664 23798
rect 11612 23734 11664 23740
rect 11716 23610 11744 24806
rect 11796 24676 11848 24682
rect 11796 24618 11848 24624
rect 11808 23714 11836 24618
rect 12176 24614 12204 26318
rect 14292 26042 14320 26998
rect 14568 26586 14596 27066
rect 14556 26580 14608 26586
rect 14556 26522 14608 26528
rect 14752 26450 14780 27406
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14844 25906 14872 27474
rect 14936 27062 14964 27542
rect 15672 27402 15700 29106
rect 15856 28762 15884 29174
rect 15844 28756 15896 28762
rect 15844 28698 15896 28704
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15764 28150 15792 28426
rect 15752 28144 15804 28150
rect 15752 28086 15804 28092
rect 15948 28082 15976 29446
rect 16040 29238 16068 31418
rect 16120 31204 16172 31210
rect 16120 31146 16172 31152
rect 16132 29578 16160 31146
rect 16224 30818 16252 31606
rect 16408 31482 16436 33918
rect 16500 33658 16528 36110
rect 16856 34944 16908 34950
rect 16856 34886 16908 34892
rect 16764 34468 16816 34474
rect 16764 34410 16816 34416
rect 16488 33652 16540 33658
rect 16488 33594 16540 33600
rect 16776 33318 16804 34410
rect 16764 33312 16816 33318
rect 16764 33254 16816 33260
rect 16868 32858 16896 34886
rect 16960 33930 16988 36518
rect 17052 36378 17080 36654
rect 17144 36582 17172 36722
rect 18064 36718 18092 39200
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18510 36816 18566 36825
rect 18510 36751 18566 36760
rect 17868 36712 17920 36718
rect 17868 36654 17920 36660
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 17132 36576 17184 36582
rect 17132 36518 17184 36524
rect 17880 36378 17908 36654
rect 17040 36372 17092 36378
rect 17040 36314 17092 36320
rect 17868 36372 17920 36378
rect 17868 36314 17920 36320
rect 18524 36310 18552 36751
rect 18512 36304 18564 36310
rect 18512 36246 18564 36252
rect 18524 36174 18552 36246
rect 18708 36242 18736 37198
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 17776 36168 17828 36174
rect 17776 36110 17828 36116
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 17684 35624 17736 35630
rect 17684 35566 17736 35572
rect 17040 35488 17092 35494
rect 17040 35430 17092 35436
rect 17052 35018 17080 35430
rect 17696 35290 17724 35566
rect 17684 35284 17736 35290
rect 17684 35226 17736 35232
rect 17040 35012 17092 35018
rect 17040 34954 17092 34960
rect 17408 35012 17460 35018
rect 17408 34954 17460 34960
rect 17052 34134 17080 34954
rect 17420 34746 17448 34954
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 17408 34604 17460 34610
rect 17408 34546 17460 34552
rect 17040 34128 17092 34134
rect 17040 34070 17092 34076
rect 16948 33924 17000 33930
rect 16948 33866 17000 33872
rect 17052 33658 17080 34070
rect 17040 33652 17092 33658
rect 17040 33594 17092 33600
rect 17420 33590 17448 34546
rect 17408 33584 17460 33590
rect 17408 33526 17460 33532
rect 16868 32842 17080 32858
rect 16868 32836 17092 32842
rect 16868 32830 17040 32836
rect 16488 32768 16540 32774
rect 16488 32710 16540 32716
rect 16500 32502 16528 32710
rect 16488 32496 16540 32502
rect 16488 32438 16540 32444
rect 16868 32366 16896 32830
rect 17040 32778 17092 32784
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 16856 32360 16908 32366
rect 16856 32302 16908 32308
rect 16764 32292 16816 32298
rect 16764 32234 16816 32240
rect 16776 32026 16804 32234
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 17236 31958 17264 32370
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 16396 31476 16448 31482
rect 16396 31418 16448 31424
rect 16500 31414 16528 31758
rect 16488 31408 16540 31414
rect 16488 31350 16540 31356
rect 16396 31340 16448 31346
rect 16396 31282 16448 31288
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16224 30790 16344 30818
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 16028 29232 16080 29238
rect 16028 29174 16080 29180
rect 16212 29164 16264 29170
rect 16212 29106 16264 29112
rect 16120 29028 16172 29034
rect 16120 28970 16172 28976
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 16132 27538 16160 28970
rect 16120 27532 16172 27538
rect 16120 27474 16172 27480
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 14924 27056 14976 27062
rect 14924 26998 14976 27004
rect 15672 26994 15700 27338
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15476 26784 15528 26790
rect 15476 26726 15528 26732
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 15384 26580 15436 26586
rect 15384 26522 15436 26528
rect 15292 26240 15344 26246
rect 15292 26182 15344 26188
rect 15304 25974 15332 26182
rect 15292 25968 15344 25974
rect 15292 25910 15344 25916
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 13096 25294 13124 25638
rect 15016 25492 15068 25498
rect 15016 25434 15068 25440
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 12268 24750 12296 25230
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12360 24818 12388 25162
rect 12452 24886 12480 25230
rect 14740 25220 14792 25226
rect 14740 25162 14792 25168
rect 14752 24954 14780 25162
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 12440 24880 12492 24886
rect 12440 24822 12492 24828
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 12164 24608 12216 24614
rect 12360 24562 12388 24754
rect 12164 24550 12216 24556
rect 12268 24534 12388 24562
rect 12268 24206 12296 24534
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 12164 24064 12216 24070
rect 12164 24006 12216 24012
rect 11900 23866 11928 24006
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 11900 23746 11928 23802
rect 11900 23730 12020 23746
rect 12176 23730 12204 24006
rect 11900 23724 12032 23730
rect 11900 23718 11980 23724
rect 11796 23708 11848 23714
rect 11980 23666 12032 23672
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 11796 23650 11848 23656
rect 11716 23582 11836 23610
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11440 22710 11468 22918
rect 11428 22704 11480 22710
rect 11428 22646 11480 22652
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11152 22500 11204 22506
rect 11152 22442 11204 22448
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 11164 21146 11192 22442
rect 11256 22030 11284 22510
rect 11336 22160 11388 22166
rect 11334 22128 11336 22137
rect 11388 22128 11390 22137
rect 11334 22063 11390 22072
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11164 21010 11192 21082
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10980 20534 11008 20878
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10980 19802 11008 20334
rect 11060 19848 11112 19854
rect 10980 19796 11060 19802
rect 10980 19790 11112 19796
rect 10980 19774 11100 19790
rect 10980 17066 11008 19774
rect 11164 19718 11192 20470
rect 11256 20398 11284 21966
rect 11348 20874 11376 21966
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11532 20602 11560 21966
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11624 21554 11652 21830
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11164 19242 11192 19654
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11624 18426 11652 19314
rect 11808 19174 11836 23582
rect 11888 23588 11940 23594
rect 12072 23588 12124 23594
rect 11940 23548 12072 23576
rect 11888 23530 11940 23536
rect 12072 23530 12124 23536
rect 12176 23202 12204 23666
rect 11992 23186 12204 23202
rect 11980 23180 12204 23186
rect 12032 23174 12204 23180
rect 11980 23122 12032 23128
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11900 22098 11928 22986
rect 12176 22982 12204 23174
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11992 22166 12020 22714
rect 12176 22642 12204 22918
rect 12268 22778 12296 24142
rect 12452 24138 12480 24822
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 12440 24132 12492 24138
rect 12440 24074 12492 24080
rect 12452 23474 12480 24074
rect 13648 23866 13676 24754
rect 13740 24342 13768 24754
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12532 23588 12584 23594
rect 12532 23530 12584 23536
rect 12360 23446 12480 23474
rect 12360 23322 12388 23446
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12360 23118 12388 23258
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12544 22778 12572 23530
rect 12912 23322 12940 23666
rect 13176 23520 13228 23526
rect 13228 23480 13308 23508
rect 13176 23462 13228 23468
rect 12900 23316 12952 23322
rect 12900 23258 12952 23264
rect 13280 23118 13308 23480
rect 13372 23118 13400 23802
rect 14108 23594 14136 24346
rect 14096 23588 14148 23594
rect 14096 23530 14148 23536
rect 14108 23118 14136 23530
rect 14200 23186 14228 24550
rect 14280 24336 14332 24342
rect 14280 24278 14332 24284
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13188 22778 13216 22986
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 13176 22772 13228 22778
rect 13176 22714 13228 22720
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12716 22568 12768 22574
rect 12768 22528 12848 22556
rect 12716 22510 12768 22516
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11900 21690 11928 22034
rect 12360 22030 12388 22374
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 12820 21554 12848 22528
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12820 20874 12848 21490
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11992 20058 12020 20402
rect 12452 20398 12480 20742
rect 12912 20534 12940 20810
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 13096 19922 13124 22034
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 13188 19854 13216 21422
rect 13372 20534 13400 23054
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13648 22030 13676 22646
rect 13832 22642 13860 23054
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 14016 22642 14044 22986
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 14004 22636 14056 22642
rect 14004 22578 14056 22584
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13648 21554 13676 21966
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13832 21146 13860 21286
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 14016 21010 14044 21626
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14004 21004 14056 21010
rect 14004 20946 14056 20952
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 11886 19544 11942 19553
rect 11886 19479 11942 19488
rect 11900 19378 11928 19479
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 13096 19174 13124 19722
rect 13372 19718 13400 19994
rect 13556 19786 13584 20810
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13648 20505 13676 20538
rect 13634 20496 13690 20505
rect 14016 20466 14044 20742
rect 13634 20431 13690 20440
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 14108 19922 14136 21490
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11256 17882 11284 18158
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11256 17678 11284 17818
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11256 17202 11284 17614
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10980 15706 11008 16050
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11440 15502 11468 18022
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11532 17542 11560 17614
rect 11624 17610 11652 18226
rect 11808 18222 11836 18702
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11624 17202 11652 17546
rect 11808 17542 11836 18158
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11624 16674 11652 17138
rect 11624 16658 11744 16674
rect 11624 16652 11756 16658
rect 11624 16646 11704 16652
rect 11704 16594 11756 16600
rect 11900 15502 11928 18770
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 16726 12020 18566
rect 12176 18154 12204 18702
rect 12268 18222 12296 18702
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12820 18154 12848 19110
rect 13096 18766 13124 19110
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 13360 18760 13412 18766
rect 13464 18748 13492 19654
rect 13740 19514 13768 19858
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13412 18720 13492 18748
rect 13360 18702 13412 18708
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13188 18204 13216 18566
rect 13280 18358 13308 18566
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13268 18216 13320 18222
rect 13188 18176 13268 18204
rect 13268 18158 13320 18164
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12176 17678 12204 18090
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17202 13032 17614
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11992 16522 12020 16662
rect 12636 16590 12664 16934
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 12912 16250 12940 17002
rect 13096 16726 13124 17138
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 12636 15434 12664 16118
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15502 12756 15846
rect 13096 15706 13124 16662
rect 13280 16658 13308 18158
rect 13372 17678 13400 18702
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13464 17134 13492 18294
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13740 16998 13768 19450
rect 13832 18290 13860 19654
rect 13910 19408 13966 19417
rect 14200 19378 14228 22170
rect 13910 19343 13966 19352
rect 14188 19372 14240 19378
rect 13924 18902 13952 19343
rect 14188 19314 14240 19320
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13924 17610 13952 18158
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 14016 16402 14044 17206
rect 14188 16448 14240 16454
rect 14016 16396 14188 16402
rect 14016 16390 14240 16396
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12544 14618 12572 15370
rect 12636 15094 12664 15370
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12728 13938 12756 14894
rect 13188 14414 13216 16390
rect 13924 16114 13952 16390
rect 14016 16374 14228 16390
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13648 14890 13676 15642
rect 13912 15632 13964 15638
rect 13912 15574 13964 15580
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 13832 13870 13860 14962
rect 13924 13938 13952 15574
rect 14016 15094 14044 16374
rect 14200 16250 14228 16374
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 12918 13860 13806
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 10520 6886 10640 6914
rect 10704 12406 10916 12434
rect 10704 6914 10732 12406
rect 13924 11898 13952 13874
rect 14016 13258 14044 14010
rect 14200 13870 14228 14214
rect 14292 14006 14320 24278
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14384 23497 14412 24074
rect 14370 23488 14426 23497
rect 14370 23423 14426 23432
rect 14476 22710 14504 24618
rect 14936 24410 14964 24754
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14660 23118 14688 23734
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14384 19417 14412 22578
rect 14476 22166 14504 22646
rect 14464 22160 14516 22166
rect 14464 22102 14516 22108
rect 14568 21418 14596 22918
rect 14660 22234 14688 23054
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14476 20534 14504 21286
rect 14844 21146 14872 21830
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14660 20602 14688 20810
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14568 19514 14596 19858
rect 14660 19854 14688 19994
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14370 19408 14426 19417
rect 14370 19343 14426 19352
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14568 18970 14596 19314
rect 14660 19310 14688 19790
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14752 17746 14780 20878
rect 14844 20398 14872 21082
rect 14924 20868 14976 20874
rect 14924 20810 14976 20816
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14936 20330 14964 20810
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 15028 19553 15056 25434
rect 15120 25362 15148 25842
rect 15396 25838 15424 26522
rect 15488 26450 15516 26726
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15948 26382 15976 26726
rect 16132 26450 16160 27474
rect 16224 27470 16252 29106
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 16224 26994 16252 27270
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 15476 26308 15528 26314
rect 15476 26250 15528 26256
rect 15488 25974 15516 26250
rect 15580 26042 15608 26318
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15476 25968 15528 25974
rect 15476 25910 15528 25916
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15384 25832 15436 25838
rect 15384 25774 15436 25780
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 15856 25294 15884 25842
rect 16224 25838 16252 26930
rect 16212 25832 16264 25838
rect 16212 25774 16264 25780
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15488 24954 15516 25094
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15488 24274 15516 24890
rect 15764 24750 15792 25094
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15580 24410 15608 24686
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15304 22438 15332 23666
rect 15488 23186 15516 24210
rect 15580 24070 15608 24346
rect 15764 24138 15792 24686
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 24138 16160 24550
rect 15752 24132 15804 24138
rect 15752 24074 15804 24080
rect 16120 24132 16172 24138
rect 16120 24074 16172 24080
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15580 23066 15608 24006
rect 15488 23050 15608 23066
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15476 23044 15608 23050
rect 15528 23038 15608 23044
rect 15476 22986 15528 22992
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 22137 15332 22374
rect 15290 22128 15346 22137
rect 15290 22063 15346 22072
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15120 20534 15148 21422
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 15120 19825 15148 20266
rect 15212 20058 15240 20402
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15106 19816 15162 19825
rect 15106 19751 15162 19760
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15014 19544 15070 19553
rect 15014 19479 15070 19488
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 17338 14596 17614
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14476 15162 14504 16458
rect 14752 16182 14780 17682
rect 14844 17066 14872 19314
rect 14924 18216 14976 18222
rect 15028 18204 15056 19479
rect 15120 19378 15148 19654
rect 15212 19446 15240 19722
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15212 18902 15240 19382
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 14976 18176 15056 18204
rect 14924 18158 14976 18164
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15212 17338 15240 17546
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15304 17270 15332 22063
rect 15488 22030 15516 22986
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15672 22642 15700 22918
rect 15764 22710 15792 23054
rect 16224 22710 16252 25162
rect 16316 24342 16344 30790
rect 16408 29646 16436 31282
rect 16488 30320 16540 30326
rect 16488 30262 16540 30268
rect 16396 29640 16448 29646
rect 16396 29582 16448 29588
rect 16408 27470 16436 29582
rect 16500 29170 16528 30262
rect 16488 29164 16540 29170
rect 16488 29106 16540 29112
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16592 26926 16620 31282
rect 16672 30864 16724 30870
rect 16672 30806 16724 30812
rect 16684 28422 16712 30806
rect 16762 30560 16818 30569
rect 16762 30495 16818 30504
rect 16776 30190 16804 30495
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16592 26518 16620 26862
rect 16580 26512 16632 26518
rect 16580 26454 16632 26460
rect 16396 25968 16448 25974
rect 16580 25968 16632 25974
rect 16448 25928 16580 25956
rect 16396 25910 16448 25916
rect 16580 25910 16632 25916
rect 16684 25906 16712 28018
rect 16776 27674 16804 28494
rect 16764 27668 16816 27674
rect 16764 27610 16816 27616
rect 16868 27606 16896 31826
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 17052 30054 17080 30670
rect 17132 30660 17184 30666
rect 17132 30602 17184 30608
rect 17144 30054 17172 30602
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17236 29646 17264 31894
rect 17420 31346 17448 33526
rect 17592 33448 17644 33454
rect 17592 33390 17644 33396
rect 17408 31340 17460 31346
rect 17408 31282 17460 31288
rect 17604 30734 17632 33390
rect 17684 31816 17736 31822
rect 17684 31758 17736 31764
rect 17696 31482 17724 31758
rect 17684 31476 17736 31482
rect 17684 31418 17736 31424
rect 17592 30728 17644 30734
rect 17592 30670 17644 30676
rect 17316 30320 17368 30326
rect 17316 30262 17368 30268
rect 17224 29640 17276 29646
rect 17224 29582 17276 29588
rect 17328 29510 17356 30262
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 28150 16988 28358
rect 17328 28218 17356 29446
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17420 28626 17448 29106
rect 17408 28620 17460 28626
rect 17408 28562 17460 28568
rect 17684 28620 17736 28626
rect 17684 28562 17736 28568
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 16948 28144 17000 28150
rect 16948 28086 17000 28092
rect 16948 28008 17000 28014
rect 16948 27950 17000 27956
rect 16856 27600 16908 27606
rect 16856 27542 16908 27548
rect 16960 26994 16988 27950
rect 17420 27674 17448 28562
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 17512 28014 17540 28494
rect 17696 28218 17724 28562
rect 17684 28212 17736 28218
rect 17684 28154 17736 28160
rect 17500 28008 17552 28014
rect 17500 27950 17552 27956
rect 17408 27668 17460 27674
rect 17408 27610 17460 27616
rect 17420 27470 17448 27610
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16960 26382 16988 26930
rect 17512 26858 17540 27950
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 17408 25968 17460 25974
rect 17408 25910 17460 25916
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24886 16620 25094
rect 16580 24880 16632 24886
rect 16580 24822 16632 24828
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 16592 23798 16620 24822
rect 16684 24206 16712 25842
rect 17420 25498 17448 25910
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 17040 25220 17092 25226
rect 17040 25162 17092 25168
rect 17052 24818 17080 25162
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17328 23798 17356 24142
rect 17788 24070 17816 36110
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 18144 35216 18196 35222
rect 18144 35158 18196 35164
rect 18156 35018 18184 35158
rect 18340 35154 18368 35430
rect 19352 35290 19380 35634
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 18340 35018 18368 35090
rect 19444 35086 19472 36518
rect 19996 36242 20024 39200
rect 20640 37330 20668 39200
rect 20628 37324 20680 37330
rect 20628 37266 20680 37272
rect 20076 37188 20128 37194
rect 20076 37130 20128 37136
rect 20088 36378 20116 37130
rect 21284 36854 21312 39200
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 21732 37120 21784 37126
rect 21732 37062 21784 37068
rect 21272 36848 21324 36854
rect 21272 36790 21324 36796
rect 21180 36780 21232 36786
rect 21180 36722 21232 36728
rect 20076 36372 20128 36378
rect 20076 36314 20128 36320
rect 19984 36236 20036 36242
rect 19984 36178 20036 36184
rect 21192 36174 21220 36722
rect 21640 36576 21692 36582
rect 21640 36518 21692 36524
rect 21180 36168 21232 36174
rect 21180 36110 21232 36116
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19522 35728 19578 35737
rect 19522 35663 19524 35672
rect 19576 35663 19578 35672
rect 20260 35692 20312 35698
rect 19524 35634 19576 35640
rect 20260 35634 20312 35640
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 20168 35080 20220 35086
rect 20168 35022 20220 35028
rect 18144 35012 18196 35018
rect 18144 34954 18196 34960
rect 18328 35012 18380 35018
rect 18328 34954 18380 34960
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 17868 34400 17920 34406
rect 17868 34342 17920 34348
rect 18512 34400 18564 34406
rect 18512 34342 18564 34348
rect 17880 34202 17908 34342
rect 17868 34196 17920 34202
rect 17868 34138 17920 34144
rect 18524 33998 18552 34342
rect 18604 34060 18656 34066
rect 18604 34002 18656 34008
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18248 33658 18276 33934
rect 18236 33652 18288 33658
rect 18236 33594 18288 33600
rect 18420 33584 18472 33590
rect 18420 33526 18472 33532
rect 18432 33114 18460 33526
rect 18616 33318 18644 34002
rect 18696 33448 18748 33454
rect 18696 33390 18748 33396
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 18420 33108 18472 33114
rect 18420 33050 18472 33056
rect 18236 32972 18288 32978
rect 18236 32914 18288 32920
rect 18052 32020 18104 32026
rect 18052 31962 18104 31968
rect 17868 31816 17920 31822
rect 17868 31758 17920 31764
rect 17880 30870 17908 31758
rect 18064 31346 18092 31962
rect 18144 31680 18196 31686
rect 18144 31622 18196 31628
rect 18156 31482 18184 31622
rect 18144 31476 18196 31482
rect 18144 31418 18196 31424
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 17960 30932 18012 30938
rect 17960 30874 18012 30880
rect 17868 30864 17920 30870
rect 17868 30806 17920 30812
rect 17972 29646 18000 30874
rect 18064 30734 18092 31282
rect 18156 30802 18184 31282
rect 18144 30796 18196 30802
rect 18144 30738 18196 30744
rect 18052 30728 18104 30734
rect 18052 30670 18104 30676
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 18064 29306 18092 30194
rect 18156 30190 18184 30738
rect 18144 30184 18196 30190
rect 18144 30126 18196 30132
rect 18248 30122 18276 32914
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 18236 30116 18288 30122
rect 18236 30058 18288 30064
rect 18340 29714 18368 32710
rect 18432 31414 18460 32846
rect 18616 32842 18644 33254
rect 18604 32836 18656 32842
rect 18604 32778 18656 32784
rect 18708 32434 18736 33390
rect 18696 32428 18748 32434
rect 18696 32370 18748 32376
rect 18892 32230 18920 34478
rect 18984 33862 19012 34546
rect 19984 34400 20036 34406
rect 19984 34342 20036 34348
rect 19996 33930 20024 34342
rect 19340 33924 19392 33930
rect 19340 33866 19392 33872
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 18972 33856 19024 33862
rect 18972 33798 19024 33804
rect 18984 33454 19012 33798
rect 18972 33448 19024 33454
rect 18972 33390 19024 33396
rect 18984 32910 19012 33390
rect 18972 32904 19024 32910
rect 18972 32846 19024 32852
rect 19156 32904 19208 32910
rect 19156 32846 19208 32852
rect 19168 32434 19196 32846
rect 19248 32564 19300 32570
rect 19248 32506 19300 32512
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19064 32360 19116 32366
rect 19064 32302 19116 32308
rect 18696 32224 18748 32230
rect 18696 32166 18748 32172
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18512 31748 18564 31754
rect 18512 31690 18564 31696
rect 18420 31408 18472 31414
rect 18420 31350 18472 31356
rect 18524 31346 18552 31690
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18708 31278 18736 32166
rect 18972 31884 19024 31890
rect 18972 31826 19024 31832
rect 18788 31748 18840 31754
rect 18788 31690 18840 31696
rect 18800 31346 18828 31690
rect 18984 31346 19012 31826
rect 19076 31482 19104 32302
rect 19260 31890 19288 32506
rect 19352 32366 19380 33866
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19524 33448 19576 33454
rect 19524 33390 19576 33396
rect 19536 32910 19564 33390
rect 19524 32904 19576 32910
rect 19444 32852 19524 32858
rect 19444 32846 19576 32852
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 19444 32830 19564 32846
rect 19444 32502 19472 32830
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19248 31884 19300 31890
rect 19248 31826 19300 31832
rect 19064 31476 19116 31482
rect 19064 31418 19116 31424
rect 19076 31346 19104 31418
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18972 31340 19024 31346
rect 18972 31282 19024 31288
rect 19064 31340 19116 31346
rect 19064 31282 19116 31288
rect 18420 31272 18472 31278
rect 18420 31214 18472 31220
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18432 30258 18460 31214
rect 19156 30796 19208 30802
rect 19156 30738 19208 30744
rect 19248 30796 19300 30802
rect 19248 30738 19300 30744
rect 19168 30258 19196 30738
rect 18420 30252 18472 30258
rect 18420 30194 18472 30200
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 19156 30252 19208 30258
rect 19156 30194 19208 30200
rect 18512 30184 18564 30190
rect 18512 30126 18564 30132
rect 18328 29708 18380 29714
rect 18328 29650 18380 29656
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18052 29300 18104 29306
rect 18052 29242 18104 29248
rect 18156 27606 18184 29582
rect 18328 29164 18380 29170
rect 18328 29106 18380 29112
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 18052 26784 18104 26790
rect 18052 26726 18104 26732
rect 18064 26586 18092 26726
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 17972 25294 18000 26182
rect 18248 25702 18276 28086
rect 18340 27470 18368 29106
rect 18524 29034 18552 30126
rect 18616 29306 18644 30194
rect 19260 30190 19288 30738
rect 19352 30258 19380 32166
rect 19432 31748 19484 31754
rect 19432 31690 19484 31696
rect 19444 31482 19472 31690
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 19996 30938 20024 31282
rect 19984 30932 20036 30938
rect 19984 30874 20036 30880
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19444 30394 19472 30670
rect 19984 30660 20036 30666
rect 19984 30602 20036 30608
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19996 30394 20024 30602
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19984 30388 20036 30394
rect 19984 30330 20036 30336
rect 20088 30258 20116 32846
rect 20180 31346 20208 35022
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19616 30252 19668 30258
rect 19616 30194 19668 30200
rect 20076 30252 20128 30258
rect 20076 30194 20128 30200
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 19248 30184 19300 30190
rect 19248 30126 19300 30132
rect 19260 30054 19288 30126
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 19352 29646 19380 30194
rect 19628 29646 19656 30194
rect 20180 29714 20208 30194
rect 20168 29708 20220 29714
rect 20168 29650 20220 29656
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19616 29640 19668 29646
rect 19616 29582 19668 29588
rect 18604 29300 18656 29306
rect 18604 29242 18656 29248
rect 18512 29028 18564 29034
rect 18512 28970 18564 28976
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 28626 18460 28902
rect 18420 28620 18472 28626
rect 18420 28562 18472 28568
rect 18432 28490 18460 28562
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 18432 27470 18460 28426
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 18340 26382 18368 26726
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17880 23798 17908 24550
rect 18340 24410 18368 25978
rect 18432 25294 18460 27066
rect 18524 26450 18552 28970
rect 18708 28694 18736 29582
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19248 29504 19300 29510
rect 19248 29446 19300 29452
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 18696 28688 18748 28694
rect 18696 28630 18748 28636
rect 18972 28552 19024 28558
rect 18972 28494 19024 28500
rect 18880 27872 18932 27878
rect 18880 27814 18932 27820
rect 18604 27532 18656 27538
rect 18604 27474 18656 27480
rect 18512 26444 18564 26450
rect 18512 26386 18564 26392
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18524 24750 18552 26386
rect 18616 26042 18644 27474
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18708 27130 18736 27270
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 18800 26790 18828 26930
rect 18892 26858 18920 27814
rect 18984 27130 19012 28494
rect 19076 27334 19104 29242
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 18972 27124 19024 27130
rect 18972 27066 19024 27072
rect 19076 26994 19104 27270
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 19076 26858 19104 26930
rect 18880 26852 18932 26858
rect 18880 26794 18932 26800
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18892 26382 18920 26794
rect 19076 26518 19104 26794
rect 19064 26512 19116 26518
rect 19064 26454 19116 26460
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 19168 25242 19196 29446
rect 19260 29170 19288 29446
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19260 28558 19288 29106
rect 19524 29028 19576 29034
rect 19524 28970 19576 28976
rect 19536 28762 19564 28970
rect 19524 28756 19576 28762
rect 19524 28698 19576 28704
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 19260 27674 19288 28018
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 19248 27668 19300 27674
rect 19248 27610 19300 27616
rect 19444 27470 19472 27882
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19444 25702 19472 27406
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 19812 26450 19840 26862
rect 19800 26444 19852 26450
rect 19800 26386 19852 26392
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 20272 25906 20300 35634
rect 20732 35086 20760 35634
rect 20812 35624 20864 35630
rect 20810 35592 20812 35601
rect 20864 35592 20866 35601
rect 20810 35527 20866 35536
rect 20720 35080 20772 35086
rect 20720 35022 20772 35028
rect 20732 34678 20760 35022
rect 20720 34672 20772 34678
rect 20720 34614 20772 34620
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20720 33584 20772 33590
rect 20720 33526 20772 33532
rect 20732 33114 20760 33526
rect 20720 33108 20772 33114
rect 20720 33050 20772 33056
rect 20824 32910 20852 34546
rect 20916 34542 20944 35974
rect 21192 35698 21220 36110
rect 21364 35760 21416 35766
rect 21364 35702 21416 35708
rect 21180 35692 21232 35698
rect 21180 35634 21232 35640
rect 20996 35556 21048 35562
rect 20996 35498 21048 35504
rect 20904 34536 20956 34542
rect 20904 34478 20956 34484
rect 21008 34202 21036 35498
rect 21376 35018 21404 35702
rect 21364 35012 21416 35018
rect 21364 34954 21416 34960
rect 20996 34196 21048 34202
rect 20996 34138 21048 34144
rect 20996 33992 21048 33998
rect 20996 33934 21048 33940
rect 21008 33590 21036 33934
rect 20996 33584 21048 33590
rect 20996 33526 21048 33532
rect 20904 33448 20956 33454
rect 20904 33390 20956 33396
rect 20916 33046 20944 33390
rect 20904 33040 20956 33046
rect 20904 32982 20956 32988
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20628 31816 20680 31822
rect 20628 31758 20680 31764
rect 20640 31482 20668 31758
rect 20824 31754 20852 32846
rect 21008 32570 21036 33526
rect 20996 32564 21048 32570
rect 20996 32506 21048 32512
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 21100 32026 21128 32370
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21376 31754 21404 34954
rect 21548 34536 21600 34542
rect 21548 34478 21600 34484
rect 21454 33008 21510 33017
rect 21454 32943 21510 32952
rect 21468 32910 21496 32943
rect 21456 32904 21508 32910
rect 21456 32846 21508 32852
rect 20732 31726 20852 31754
rect 21192 31726 21404 31754
rect 20628 31476 20680 31482
rect 20628 31418 20680 31424
rect 20732 31346 20760 31726
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20732 30258 20760 31282
rect 20904 31272 20956 31278
rect 20904 31214 20956 31220
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20824 30326 20852 30534
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20824 29714 20852 30262
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20824 28608 20852 29650
rect 20916 29170 20944 31214
rect 20996 30660 21048 30666
rect 20996 30602 21048 30608
rect 21008 30394 21036 30602
rect 20996 30388 21048 30394
rect 20996 30330 21048 30336
rect 21088 29572 21140 29578
rect 21088 29514 21140 29520
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20904 28620 20956 28626
rect 20824 28580 20904 28608
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20640 27470 20668 28154
rect 20444 27464 20496 27470
rect 20444 27406 20496 27412
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20352 27328 20404 27334
rect 20352 27270 20404 27276
rect 20364 26314 20392 27270
rect 20456 27130 20484 27406
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 19076 25214 19196 25242
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 16580 23792 16632 23798
rect 16580 23734 16632 23740
rect 17224 23792 17276 23798
rect 17224 23734 17276 23740
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 16212 22704 16264 22710
rect 16212 22646 16264 22652
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15764 22098 15792 22646
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15856 21962 15884 22578
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15580 20806 15608 21490
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15580 20534 15608 20742
rect 15856 20602 15884 21490
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 19990 15424 20198
rect 15580 20058 15608 20470
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 15856 19854 15884 20538
rect 16132 20058 16160 22578
rect 16408 22166 16436 23122
rect 16684 22506 16712 23666
rect 16868 23322 16896 23666
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17052 23118 17080 23190
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 16396 22160 16448 22166
rect 16396 22102 16448 22108
rect 16776 22094 16804 23054
rect 17236 22982 17264 23734
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17512 23118 17540 23462
rect 19076 23322 19104 25214
rect 19156 25152 19208 25158
rect 19156 25094 19208 25100
rect 19168 24886 19196 25094
rect 19156 24880 19208 24886
rect 19156 24822 19208 24828
rect 19260 24206 19288 25230
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19260 23730 19288 24142
rect 19248 23724 19300 23730
rect 19248 23666 19300 23672
rect 19064 23316 19116 23322
rect 19064 23258 19116 23264
rect 19444 23254 19472 25434
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 20088 23866 20116 25162
rect 20168 24132 20220 24138
rect 20168 24074 20220 24080
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 16684 22066 16804 22094
rect 16684 22030 16712 22066
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16408 21486 16436 21898
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16408 21010 16436 21422
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15580 18766 15608 19110
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15396 17202 15424 18566
rect 15764 18290 15792 19110
rect 15856 18970 15884 19790
rect 16040 19242 16068 19994
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15856 17882 15884 18906
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 15752 16720 15804 16726
rect 15752 16662 15804 16668
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14752 15638 14780 16118
rect 15764 16114 15792 16662
rect 15856 16590 15884 17478
rect 16316 17202 16344 19994
rect 16408 19446 16436 20946
rect 16592 20942 16620 21286
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16592 20534 16620 20878
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16592 19854 16620 20470
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 16408 18698 16436 19382
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16500 17610 16528 18566
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16592 18086 16620 18158
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16684 17746 16712 19926
rect 16776 19922 16804 20198
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16868 19854 16896 21354
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16762 19544 16818 19553
rect 16762 19479 16764 19488
rect 16816 19479 16818 19488
rect 16764 19450 16816 19456
rect 16960 19292 16988 22714
rect 17236 22642 17264 22918
rect 17512 22710 17540 23054
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17972 22234 18000 23054
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17960 22228 18012 22234
rect 17960 22170 18012 22176
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 19514 17080 20198
rect 17144 19786 17172 21966
rect 18064 21622 18092 22918
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18156 21622 18184 22578
rect 18248 22098 18276 23054
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22710 18920 22918
rect 18880 22704 18932 22710
rect 18880 22646 18932 22652
rect 18236 22092 18288 22098
rect 18892 22094 18920 22646
rect 19444 22574 19472 23054
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19352 22094 19380 22374
rect 18892 22066 19104 22094
rect 18236 22034 18288 22040
rect 18420 21956 18472 21962
rect 18420 21898 18472 21904
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 20534 18092 21422
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18052 20528 18104 20534
rect 17866 20496 17922 20505
rect 18052 20470 18104 20476
rect 17866 20431 17922 20440
rect 17880 20398 17908 20431
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17224 19848 17276 19854
rect 17328 19825 17356 19926
rect 17500 19848 17552 19854
rect 17224 19790 17276 19796
rect 17314 19816 17370 19825
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17236 19378 17264 19790
rect 17500 19790 17552 19796
rect 17314 19751 17370 19760
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 16868 19264 16988 19292
rect 16868 18086 16896 19264
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16960 18426 16988 18566
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17052 18222 17080 18702
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16500 16590 16528 17546
rect 16592 16590 16620 17614
rect 16684 17338 16712 17682
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16776 16590 16804 18022
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16960 16794 16988 17138
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17052 16658 17080 18158
rect 17236 18154 17264 18770
rect 17328 18698 17356 19751
rect 17512 18834 17540 19790
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17696 18766 17724 18838
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 18064 18698 18092 19110
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 17236 17678 17264 18090
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 18156 17270 18184 20742
rect 18248 20262 18276 20946
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18248 19922 18276 20198
rect 18340 20058 18368 20538
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18248 19446 18276 19858
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18340 19514 18368 19654
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18236 19440 18288 19446
rect 18432 19417 18460 21898
rect 19076 21486 19104 22066
rect 19168 22066 19380 22094
rect 19444 22094 19472 22510
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19628 22166 19656 22374
rect 19616 22160 19668 22166
rect 19616 22102 19668 22108
rect 19904 22098 19932 22646
rect 19996 22574 20024 23666
rect 20088 23118 20116 23802
rect 20180 23526 20208 24074
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20180 23118 20208 23462
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19444 22066 19564 22094
rect 19168 22030 19196 22066
rect 19156 22024 19208 22030
rect 19536 21978 19564 22066
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19156 21966 19208 21972
rect 19352 21950 19564 21978
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19260 21622 19288 21830
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19352 21554 19380 21950
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18236 19382 18288 19388
rect 18418 19408 18474 19417
rect 18418 19343 18474 19352
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18248 18086 18276 18770
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18432 17746 18460 19343
rect 18524 18834 18552 19994
rect 18616 19553 18644 21422
rect 19444 21418 19472 21830
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19996 21554 20024 22510
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18602 19544 18658 19553
rect 18602 19479 18658 19488
rect 18708 18902 18736 21286
rect 19444 21078 19472 21354
rect 20088 21146 20116 21830
rect 20272 21690 20300 25638
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20364 23662 20392 25298
rect 20640 25294 20668 27406
rect 20824 26994 20852 28580
rect 20904 28562 20956 28568
rect 21008 28490 21036 29446
rect 21100 29306 21128 29514
rect 21088 29300 21140 29306
rect 21088 29242 21140 29248
rect 21192 29186 21220 31726
rect 21100 29158 21220 29186
rect 20996 28484 21048 28490
rect 20996 28426 21048 28432
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20732 25888 20760 26726
rect 20824 26450 20852 26930
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 20812 26444 20864 26450
rect 20812 26386 20864 26392
rect 20916 25974 20944 26726
rect 20904 25968 20956 25974
rect 20904 25910 20956 25916
rect 20732 25860 20852 25888
rect 20824 25770 20852 25860
rect 20720 25764 20772 25770
rect 20720 25706 20772 25712
rect 20812 25764 20864 25770
rect 20812 25706 20864 25712
rect 20732 25294 20760 25706
rect 21008 25702 21036 26726
rect 21100 26246 21128 29158
rect 21180 29028 21232 29034
rect 21180 28970 21232 28976
rect 21192 27130 21220 28970
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 21376 28218 21404 28494
rect 21364 28212 21416 28218
rect 21364 28154 21416 28160
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 21180 27124 21232 27130
rect 21180 27066 21232 27072
rect 21272 27056 21324 27062
rect 21272 26998 21324 27004
rect 21284 26586 21312 26998
rect 21272 26580 21324 26586
rect 21272 26522 21324 26528
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21284 25974 21312 26522
rect 21272 25968 21324 25974
rect 21272 25910 21324 25916
rect 21468 25770 21496 27814
rect 21456 25764 21508 25770
rect 21456 25706 21508 25712
rect 20996 25696 21048 25702
rect 20916 25644 20996 25650
rect 20916 25638 21048 25644
rect 20916 25622 21036 25638
rect 20916 25430 20944 25622
rect 21468 25498 21496 25706
rect 21456 25492 21508 25498
rect 21456 25434 21508 25440
rect 20904 25424 20956 25430
rect 20904 25366 20956 25372
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20732 24886 20760 25230
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20640 23730 20668 24074
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 19432 21072 19484 21078
rect 19432 21014 19484 21020
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19168 19786 19196 20402
rect 19352 20074 19380 20878
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19996 20602 20024 20878
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19260 20046 19380 20074
rect 19156 19780 19208 19786
rect 19156 19722 19208 19728
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18800 18902 18828 19246
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18432 17270 18460 17682
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18524 17202 18552 18566
rect 18616 17882 18644 18702
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18708 17678 18736 18838
rect 18984 17678 19012 19314
rect 19168 19310 19196 19722
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19168 18630 19196 19246
rect 19260 19242 19288 20046
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19352 18358 19380 19926
rect 19444 19310 19472 20470
rect 19996 20398 20024 20538
rect 20272 20398 20300 20742
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19446 20024 20198
rect 20088 19514 20116 20334
rect 20364 20058 20392 23598
rect 20548 23186 20576 23666
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20456 21554 20484 22918
rect 20534 22536 20590 22545
rect 20640 22522 20668 23666
rect 20590 22494 20668 22522
rect 20534 22471 20590 22480
rect 20548 22234 20576 22471
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20916 21622 20944 25366
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 21284 25265 21312 25298
rect 21270 25256 21326 25265
rect 21270 25191 21326 25200
rect 21284 24954 21312 25191
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 17882 19288 18226
rect 19352 17882 19380 18294
rect 19444 18290 19472 19246
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 20088 18426 20116 19450
rect 20352 18964 20404 18970
rect 20456 18952 20484 20810
rect 20404 18924 20484 18952
rect 20352 18906 20404 18912
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18984 17338 19012 17614
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16764 16584 16816 16590
rect 17972 16572 18000 17138
rect 19444 17134 19472 18226
rect 20364 18086 20392 18226
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20364 17746 20392 18022
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19246 16688 19302 16697
rect 19246 16623 19302 16632
rect 16764 16526 16816 16532
rect 17880 16544 18000 16572
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15120 15162 15148 15370
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14476 14006 14504 14758
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14568 13870 14596 14486
rect 15212 14074 15240 14962
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14016 12170 14044 12582
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13096 9586 13124 11834
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14200 11354 14228 11630
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14292 10810 14320 11698
rect 14384 11150 14412 12038
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9654 14136 9862
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13464 9178 13492 9454
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8634 13584 8910
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 10704 6886 10916 6914
rect 10520 4622 10548 6886
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 9140 2378 9168 3334
rect 9232 3126 9260 3878
rect 10612 3602 10640 3878
rect 10796 3602 10824 4626
rect 10888 4146 10916 6886
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 9692 800 9720 2926
rect 10980 800 11008 3606
rect 11256 3602 11284 3878
rect 11440 3602 11468 4422
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 13372 2446 13400 3674
rect 13832 3058 13860 3878
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14292 3058 14320 3538
rect 14568 3534 14596 13806
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13530 15516 13670
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 11830 15240 12786
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15212 10674 15240 11766
rect 15580 11762 15608 14962
rect 15764 14958 15792 16050
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 15856 15434 15884 15846
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 16684 14958 16712 15846
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15672 13530 15700 14350
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10810 15332 11086
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15212 10062 15240 10610
rect 15396 10062 15424 10610
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 8906 14872 9862
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15212 8090 15240 8434
rect 15396 8430 15424 9998
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15488 9178 15516 9386
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15580 9042 15608 10406
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15672 8430 15700 10542
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15396 7886 15424 8366
rect 15764 7886 15792 14350
rect 15948 13870 15976 14350
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 16592 13326 16620 14214
rect 16684 13394 16712 14894
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16580 13320 16632 13326
rect 16776 13274 16804 13806
rect 16580 13262 16632 13268
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 16684 13246 16804 13274
rect 16132 12986 16160 13194
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16684 12850 16712 13246
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16776 12850 16804 13126
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15948 11218 15976 12174
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15856 9178 15884 10542
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15948 9042 15976 11154
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7546 15792 7686
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14844 6458 14872 6666
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 15396 6322 15424 7142
rect 15948 6882 15976 8978
rect 15856 6866 15976 6882
rect 15844 6860 15976 6866
rect 15896 6854 15976 6860
rect 15844 6802 15896 6808
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15488 5914 15516 6666
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15948 5166 15976 6854
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16040 5370 16068 5646
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16132 5234 16160 11698
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16408 10810 16436 11154
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9518 16620 9998
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16592 9382 16620 9454
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16684 8634 16712 10610
rect 16776 10470 16804 12242
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 10538 16896 11494
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16776 9382 16804 10406
rect 16868 10198 16896 10474
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16960 9654 16988 12786
rect 17052 12374 17080 14350
rect 17144 12918 17172 16050
rect 17880 16046 17908 16544
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17328 14618 17356 14894
rect 17512 14618 17540 15302
rect 17696 15162 17724 15438
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17236 14006 17264 14486
rect 17512 14006 17540 14554
rect 17696 14346 17724 15098
rect 17880 14618 17908 15438
rect 17972 15094 18000 16390
rect 18156 16182 18184 16390
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18248 15706 18276 15982
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18892 15094 18920 15642
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 18880 15088 18932 15094
rect 18880 15030 18932 15036
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17880 14278 17908 14554
rect 17972 14414 18000 14894
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14618 19104 14758
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17328 13394 17356 13738
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 17052 11762 17080 12310
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17144 10742 17172 12854
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11898 17356 12038
rect 17512 11898 17540 13330
rect 17972 12306 18000 14214
rect 18064 13530 18092 14282
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18248 13258 18276 14350
rect 18524 13954 18552 14350
rect 18432 13938 18552 13954
rect 18420 13932 18552 13938
rect 18472 13926 18552 13932
rect 18696 13932 18748 13938
rect 18420 13874 18472 13880
rect 18696 13874 18748 13880
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17328 10062 17356 11290
rect 17788 11082 17816 12038
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17972 11218 18000 11834
rect 18064 11694 18092 12174
rect 18248 11898 18276 13194
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12442 18368 13126
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17788 10742 17816 11018
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16868 8906 16896 9590
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16868 8498 16896 8842
rect 17052 8498 17080 9046
rect 17236 8974 17264 9454
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17144 8498 17172 8774
rect 17420 8634 17448 9522
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16408 7546 16436 7822
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16960 7478 16988 8298
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16684 6866 16712 7278
rect 16856 7268 16908 7274
rect 16856 7210 16908 7216
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16684 5914 16712 6054
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15948 4690 15976 5102
rect 16132 4690 16160 5170
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16592 4554 16620 5510
rect 16776 4826 16804 6598
rect 16868 6390 16896 7210
rect 16960 6798 16988 7414
rect 17052 7342 17080 7822
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17052 6458 17080 6802
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 17420 5710 17448 8570
rect 17512 8498 17540 8978
rect 17604 8974 17632 10202
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17696 8514 17724 10542
rect 17972 9654 18000 11154
rect 18064 11014 18092 11630
rect 18340 11558 18368 12378
rect 18616 11898 18644 13806
rect 18708 12986 18736 13874
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18708 12306 18736 12786
rect 18800 12782 18828 14350
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18984 12900 19012 14282
rect 19076 13870 19104 14554
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19260 13734 19288 16623
rect 19352 14822 19380 16730
rect 19444 16658 19472 17070
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19812 15570 19840 15846
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19444 15026 19472 15302
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19352 14074 19380 14486
rect 19720 14482 19748 14758
rect 19904 14634 19932 14962
rect 19996 14822 20024 15302
rect 20088 15178 20116 16390
rect 20180 16250 20208 17070
rect 20260 16652 20312 16658
rect 20548 16640 20576 21286
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20718 20088 20774 20097
rect 20718 20023 20774 20032
rect 20732 19922 20760 20023
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20732 19825 20760 19858
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20824 18766 20852 20198
rect 20916 19718 20944 20878
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20916 19174 20944 19654
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20548 16612 20668 16640
rect 20260 16594 20312 16600
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20088 15150 20208 15178
rect 20272 15162 20300 16594
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 16250 20484 16390
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20180 15042 20208 15150
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20180 15014 20300 15042
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19904 14606 20024 14634
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19352 12986 19380 13738
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19064 12912 19116 12918
rect 18984 12872 19064 12900
rect 19064 12854 19116 12860
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18708 11762 18736 12242
rect 18800 12170 18828 12718
rect 19076 12481 19104 12854
rect 19062 12472 19118 12481
rect 19062 12407 19118 12416
rect 19168 12434 19196 12854
rect 19444 12850 19472 14214
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19996 13802 20024 14606
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19984 13184 20036 13190
rect 20088 13172 20116 14894
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20036 13144 20116 13172
rect 19984 13126 20036 13132
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19996 12714 20024 13126
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19168 12406 19288 12434
rect 19260 12170 19288 12406
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 11218 18644 11494
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18708 11082 18736 11698
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10810 18092 10950
rect 18708 10810 18736 11018
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18064 10266 18092 10610
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18064 9722 18092 10202
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9178 18092 9454
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17880 8906 17908 9046
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17696 8498 17908 8514
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17696 8492 17920 8498
rect 17696 8486 17868 8492
rect 17696 7478 17724 8486
rect 17868 8434 17920 8440
rect 17972 7970 18000 8910
rect 18064 8362 18092 9114
rect 18156 8974 18184 10678
rect 18800 10130 18828 12106
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17788 7942 18000 7970
rect 17788 7562 17816 7942
rect 17972 7818 18000 7942
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17880 7698 17908 7754
rect 18064 7698 18092 8298
rect 18156 8090 18184 8910
rect 18248 8634 18276 9658
rect 18340 8906 18368 9930
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18248 8362 18276 8570
rect 18616 8378 18644 9386
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18524 8350 18644 8378
rect 18524 8090 18552 8350
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18236 7744 18288 7750
rect 17880 7670 18184 7698
rect 18236 7686 18288 7692
rect 17788 7534 18000 7562
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17696 7274 17724 7414
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17972 6458 18000 7534
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17696 5914 17724 6258
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17972 5710 18000 6394
rect 18156 6390 18184 7670
rect 18248 6866 18276 7686
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18432 7206 18460 7482
rect 18524 7478 18552 8026
rect 18708 7886 18736 9590
rect 18892 9586 18920 9930
rect 18984 9586 19012 9998
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18800 8566 18828 8910
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18800 8022 18828 8502
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18892 7546 18920 8774
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18524 7342 18552 7414
rect 18984 7410 19012 9522
rect 19076 8566 19104 11766
rect 19260 11762 19288 12106
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19168 9994 19196 10610
rect 19352 10033 19380 12650
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19444 10470 19472 11630
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19720 10266 19748 10406
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19904 10146 19932 10542
rect 19996 10266 20024 11698
rect 20088 11558 20116 12174
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 20088 10198 20116 11018
rect 20076 10192 20128 10198
rect 19904 10118 20024 10146
rect 20076 10134 20128 10140
rect 19338 10024 19394 10033
rect 19156 9988 19208 9994
rect 19338 9959 19394 9968
rect 19156 9930 19208 9936
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9654 19288 9862
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18432 6798 18460 7142
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 18064 5778 18092 6258
rect 18432 6186 18460 6734
rect 18524 6322 18552 7142
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 16868 4826 16896 5646
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17144 5302 17172 5510
rect 18524 5370 18552 5646
rect 18616 5370 18644 6122
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17868 5296 17920 5302
rect 17868 5238 17920 5244
rect 17880 4826 17908 5238
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 18524 4622 18552 5306
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 18708 4146 18736 6598
rect 18800 6390 18828 6598
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18984 5710 19012 6258
rect 19168 6186 19196 9522
rect 19352 9466 19380 9959
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19260 9438 19380 9466
rect 19260 9178 19288 9438
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19352 8498 19380 9318
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19444 8566 19472 9046
rect 19904 8820 19932 9522
rect 19996 9382 20024 10118
rect 20088 9586 20116 10134
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 8974 20024 9318
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 20074 8936 20130 8945
rect 20074 8871 20130 8880
rect 20088 8838 20116 8871
rect 20076 8832 20128 8838
rect 19904 8792 20024 8820
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19352 7274 19380 7754
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19444 7313 19472 7346
rect 19430 7304 19486 7313
rect 19340 7268 19392 7274
rect 19430 7239 19486 7248
rect 19340 7210 19392 7216
rect 19156 6180 19208 6186
rect 19156 6122 19208 6128
rect 19352 5930 19380 7210
rect 19536 6712 19564 7346
rect 19996 6730 20024 8792
rect 20076 8774 20128 8780
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20088 7546 20116 8434
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20180 7410 20208 13874
rect 20272 11150 20300 15014
rect 20364 13530 20392 16050
rect 20548 15978 20576 16458
rect 20640 16182 20668 16612
rect 20732 16522 20760 17478
rect 21008 17082 21036 24006
rect 21192 23225 21220 24210
rect 21178 23216 21234 23225
rect 21178 23151 21234 23160
rect 21192 23118 21220 23151
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21192 22438 21220 23054
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 20824 17054 21036 17082
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20444 15632 20496 15638
rect 20444 15574 20496 15580
rect 20456 13938 20484 15574
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20272 8945 20300 11086
rect 20258 8936 20314 8945
rect 20258 8871 20314 8880
rect 20364 8634 20392 13262
rect 20456 11830 20484 13670
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20548 11558 20576 15302
rect 20824 15178 20852 17054
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 15502 20944 16934
rect 21100 16538 21128 21286
rect 21192 21146 21220 21422
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 17270 21220 17478
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 21100 16510 21220 16538
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21100 16114 21128 16390
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21100 15570 21128 16050
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20732 15150 20852 15178
rect 20732 14634 20760 15150
rect 20916 15094 20944 15302
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 21008 15026 21036 15098
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20640 14606 20760 14634
rect 20640 14550 20668 14606
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20732 13938 20760 14486
rect 20824 14482 20852 14962
rect 20902 14648 20958 14657
rect 20902 14583 20904 14592
rect 20956 14583 20958 14592
rect 20904 14554 20956 14560
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 21008 14362 21036 14962
rect 20916 14334 21036 14362
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20824 13870 20852 13942
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20640 13462 20668 13670
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12986 20760 13126
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20640 12102 20668 12786
rect 20916 12782 20944 14334
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 21008 13394 21036 14214
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 21100 13274 21128 13466
rect 21008 13258 21128 13274
rect 20996 13252 21128 13258
rect 21048 13246 21128 13252
rect 20996 13194 21048 13200
rect 21008 12918 21036 13194
rect 21192 12918 21220 16510
rect 20996 12912 21048 12918
rect 21180 12912 21232 12918
rect 21048 12872 21128 12900
rect 20996 12854 21048 12860
rect 21100 12782 21128 12872
rect 21180 12854 21232 12860
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20916 12238 20944 12718
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11898 20668 12038
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20456 10146 20484 11494
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20812 11008 20864 11014
rect 20640 10968 20812 10996
rect 20640 10606 20668 10968
rect 20812 10950 20864 10956
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20548 10266 20576 10406
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20456 10118 20576 10146
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20364 7342 20392 8570
rect 20352 7336 20404 7342
rect 20272 7296 20352 7324
rect 19260 5902 19380 5930
rect 19444 6684 19564 6712
rect 19984 6724 20036 6730
rect 19444 5914 19472 6684
rect 19984 6666 20036 6672
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19996 6390 20024 6666
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19432 5908 19484 5914
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 19260 5574 19288 5902
rect 19432 5850 19484 5856
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19352 5302 19380 5714
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19904 5658 19932 6054
rect 20272 5914 20300 7296
rect 20352 7278 20404 7284
rect 20352 6384 20404 6390
rect 20352 6326 20404 6332
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19444 5030 19472 5646
rect 19904 5630 20024 5658
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19996 5166 20024 5630
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19444 4690 19472 4966
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19996 4282 20024 4490
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 20088 4010 20116 5578
rect 20364 5370 20392 6326
rect 20456 6254 20484 9930
rect 20548 8498 20576 10118
rect 20824 9722 20852 10610
rect 20916 10538 20944 11086
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 21008 10266 21036 10542
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20916 9518 20944 9658
rect 20904 9512 20956 9518
rect 21100 9466 21128 12718
rect 21192 12238 21220 12854
rect 21284 12434 21312 24754
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21376 22642 21404 23054
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21376 22098 21404 22578
rect 21468 22273 21496 23258
rect 21454 22264 21510 22273
rect 21454 22199 21510 22208
rect 21364 22092 21416 22098
rect 21560 22094 21588 34478
rect 21652 24818 21680 36518
rect 21744 35834 21772 37062
rect 21732 35828 21784 35834
rect 21732 35770 21784 35776
rect 21836 35562 21864 37198
rect 22376 37188 22428 37194
rect 22376 37130 22428 37136
rect 21916 37120 21968 37126
rect 21916 37062 21968 37068
rect 21928 36718 21956 37062
rect 21916 36712 21968 36718
rect 21916 36654 21968 36660
rect 22008 36304 22060 36310
rect 22008 36246 22060 36252
rect 22020 35698 22048 36246
rect 22388 36106 22416 37130
rect 22836 37120 22888 37126
rect 22836 37062 22888 37068
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22376 36100 22428 36106
rect 22376 36042 22428 36048
rect 22388 36009 22416 36042
rect 22374 36000 22430 36009
rect 22374 35935 22430 35944
rect 22664 35698 22692 36110
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 22652 35692 22704 35698
rect 22652 35634 22704 35640
rect 21824 35556 21876 35562
rect 21824 35498 21876 35504
rect 21916 34740 21968 34746
rect 21916 34682 21968 34688
rect 21928 34066 21956 34682
rect 21916 34060 21968 34066
rect 21916 34002 21968 34008
rect 21732 32836 21784 32842
rect 21732 32778 21784 32784
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21744 22094 21772 32778
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21824 29504 21876 29510
rect 21824 29446 21876 29452
rect 21836 29170 21864 29446
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 21928 27878 21956 31758
rect 22020 31210 22048 35634
rect 22848 35630 22876 37062
rect 23124 36922 23152 37198
rect 23112 36916 23164 36922
rect 23112 36858 23164 36864
rect 22836 35624 22888 35630
rect 22836 35566 22888 35572
rect 22468 34604 22520 34610
rect 22468 34546 22520 34552
rect 22480 33658 22508 34546
rect 22652 33924 22704 33930
rect 22652 33866 22704 33872
rect 22468 33652 22520 33658
rect 22468 33594 22520 33600
rect 22664 33114 22692 33866
rect 22652 33108 22704 33114
rect 22652 33050 22704 33056
rect 22928 32768 22980 32774
rect 22928 32710 22980 32716
rect 22560 32496 22612 32502
rect 22560 32438 22612 32444
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22112 31822 22140 32166
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 22572 31482 22600 32438
rect 22836 31884 22888 31890
rect 22836 31826 22888 31832
rect 22848 31482 22876 31826
rect 22940 31754 22968 32710
rect 22928 31748 22980 31754
rect 22928 31690 22980 31696
rect 22560 31476 22612 31482
rect 22560 31418 22612 31424
rect 22836 31476 22888 31482
rect 22836 31418 22888 31424
rect 22008 31204 22060 31210
rect 22008 31146 22060 31152
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22192 30660 22244 30666
rect 22192 30602 22244 30608
rect 22204 30394 22232 30602
rect 22192 30388 22244 30394
rect 22192 30330 22244 30336
rect 22572 30258 22600 31078
rect 22928 30660 22980 30666
rect 22928 30602 22980 30608
rect 22940 30326 22968 30602
rect 22928 30320 22980 30326
rect 22928 30262 22980 30268
rect 22560 30252 22612 30258
rect 22560 30194 22612 30200
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22652 29572 22704 29578
rect 22652 29514 22704 29520
rect 22008 29096 22060 29102
rect 22008 29038 22060 29044
rect 22020 28218 22048 29038
rect 22664 28218 22692 29514
rect 22008 28212 22060 28218
rect 22008 28154 22060 28160
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22848 28082 22876 30126
rect 22928 28552 22980 28558
rect 22928 28494 22980 28500
rect 22940 28150 22968 28494
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 21916 27872 21968 27878
rect 21916 27814 21968 27820
rect 21916 27668 21968 27674
rect 21916 27610 21968 27616
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21836 26382 21864 27066
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 24206 21864 24754
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21928 22094 21956 27610
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22008 26308 22060 26314
rect 22008 26250 22060 26256
rect 22020 25702 22048 26250
rect 22112 26042 22140 26862
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22204 25922 22232 28018
rect 22284 27600 22336 27606
rect 22284 27542 22336 27548
rect 22296 26518 22324 27542
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 27062 22784 27270
rect 22744 27056 22796 27062
rect 22744 26998 22796 27004
rect 22284 26512 22336 26518
rect 22284 26454 22336 26460
rect 22560 26376 22612 26382
rect 22560 26318 22612 26324
rect 22112 25894 22232 25922
rect 22284 25900 22336 25906
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 22112 24750 22140 25894
rect 22284 25842 22336 25848
rect 22296 25498 22324 25842
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22572 25294 22600 26318
rect 22744 25832 22796 25838
rect 22744 25774 22796 25780
rect 22756 25294 22784 25774
rect 22848 25498 22876 28018
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22940 25294 22968 28086
rect 23124 25430 23152 36858
rect 23216 35630 23244 39200
rect 23664 37256 23716 37262
rect 23664 37198 23716 37204
rect 24124 37256 24176 37262
rect 24124 37198 24176 37204
rect 23676 36786 23704 37198
rect 24136 36786 24164 37198
rect 24504 36802 24532 39200
rect 25412 37256 25464 37262
rect 25412 37198 25464 37204
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 26148 37256 26200 37262
rect 26148 37198 26200 37204
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 24124 36780 24176 36786
rect 24504 36774 24624 36802
rect 24124 36722 24176 36728
rect 24596 36718 24624 36774
rect 24492 36712 24544 36718
rect 24492 36654 24544 36660
rect 24584 36712 24636 36718
rect 24584 36654 24636 36660
rect 24504 36378 24532 36654
rect 24492 36372 24544 36378
rect 24492 36314 24544 36320
rect 25424 36242 25452 37198
rect 25792 36922 25820 37198
rect 25964 37120 26016 37126
rect 25964 37062 26016 37068
rect 25780 36916 25832 36922
rect 25780 36858 25832 36864
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 23204 35624 23256 35630
rect 23204 35566 23256 35572
rect 24596 35290 24624 36110
rect 25044 36032 25096 36038
rect 25044 35974 25096 35980
rect 24584 35284 24636 35290
rect 24584 35226 24636 35232
rect 23664 34944 23716 34950
rect 23664 34886 23716 34892
rect 23676 34678 23704 34886
rect 23664 34672 23716 34678
rect 23664 34614 23716 34620
rect 24124 34128 24176 34134
rect 24124 34070 24176 34076
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23400 33590 23428 34002
rect 23480 33856 23532 33862
rect 23480 33798 23532 33804
rect 23388 33584 23440 33590
rect 23388 33526 23440 33532
rect 23492 33454 23520 33798
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 23480 33448 23532 33454
rect 23480 33390 23532 33396
rect 23492 32910 23520 33390
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23388 32904 23440 32910
rect 23388 32846 23440 32852
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23400 31822 23428 32846
rect 23584 32774 23612 33254
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 24044 32502 24072 33458
rect 24032 32496 24084 32502
rect 24032 32438 24084 32444
rect 23572 32360 23624 32366
rect 23572 32302 23624 32308
rect 23584 31890 23612 32302
rect 24136 32026 24164 34070
rect 24216 33992 24268 33998
rect 24596 33969 24624 35226
rect 24860 35148 24912 35154
rect 24860 35090 24912 35096
rect 24872 34746 24900 35090
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 25056 34678 25084 35974
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 25148 35018 25176 35430
rect 25136 35012 25188 35018
rect 25136 34954 25188 34960
rect 25228 34944 25280 34950
rect 25228 34886 25280 34892
rect 25044 34672 25096 34678
rect 25044 34614 25096 34620
rect 25044 34536 25096 34542
rect 25044 34478 25096 34484
rect 24676 33992 24728 33998
rect 24216 33934 24268 33940
rect 24582 33960 24638 33969
rect 24228 32774 24256 33934
rect 24676 33934 24728 33940
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 24582 33895 24638 33904
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 24412 33658 24440 33798
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 24688 33538 24716 33934
rect 24964 33658 24992 33934
rect 24952 33652 25004 33658
rect 24952 33594 25004 33600
rect 24596 33510 24716 33538
rect 25056 33522 25084 34478
rect 25240 34202 25268 34886
rect 25228 34196 25280 34202
rect 25228 34138 25280 34144
rect 25228 33584 25280 33590
rect 25228 33526 25280 33532
rect 25044 33516 25096 33522
rect 24596 33454 24624 33510
rect 25044 33458 25096 33464
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24860 33448 24912 33454
rect 24860 33390 24912 33396
rect 24400 33312 24452 33318
rect 24872 33300 24900 33390
rect 24400 33254 24452 33260
rect 24596 33272 24900 33300
rect 24952 33312 25004 33318
rect 24412 33046 24440 33254
rect 24596 33114 24624 33272
rect 24952 33254 25004 33260
rect 24584 33108 24636 33114
rect 24584 33050 24636 33056
rect 24400 33040 24452 33046
rect 24400 32982 24452 32988
rect 24308 32836 24360 32842
rect 24308 32778 24360 32784
rect 24216 32768 24268 32774
rect 24216 32710 24268 32716
rect 24228 32366 24256 32710
rect 24320 32366 24348 32778
rect 24216 32360 24268 32366
rect 24216 32302 24268 32308
rect 24308 32360 24360 32366
rect 24308 32302 24360 32308
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23400 31414 23428 31758
rect 24228 31482 24256 32302
rect 24320 31822 24348 32302
rect 24412 32026 24440 32982
rect 24492 32904 24544 32910
rect 24492 32846 24544 32852
rect 24504 32366 24532 32846
rect 24964 32774 24992 33254
rect 25056 32842 25084 33458
rect 25044 32836 25096 32842
rect 25044 32778 25096 32784
rect 24952 32768 25004 32774
rect 24952 32710 25004 32716
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24492 32360 24544 32366
rect 24492 32302 24544 32308
rect 24400 32020 24452 32026
rect 24400 31962 24452 31968
rect 24308 31816 24360 31822
rect 24308 31758 24360 31764
rect 24320 31482 24348 31758
rect 24400 31748 24452 31754
rect 24400 31690 24452 31696
rect 24216 31476 24268 31482
rect 24216 31418 24268 31424
rect 24308 31476 24360 31482
rect 24308 31418 24360 31424
rect 23388 31408 23440 31414
rect 23388 31350 23440 31356
rect 23400 30258 23428 31350
rect 24412 31278 24440 31690
rect 23664 31272 23716 31278
rect 23664 31214 23716 31220
rect 24400 31272 24452 31278
rect 24400 31214 24452 31220
rect 23676 30938 23704 31214
rect 23480 30932 23532 30938
rect 23480 30874 23532 30880
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 23400 29646 23428 30194
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23492 29306 23520 30874
rect 24400 29708 24452 29714
rect 24400 29650 24452 29656
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23492 27470 23520 29242
rect 23572 29232 23624 29238
rect 23572 29174 23624 29180
rect 23584 28626 23612 29174
rect 23572 28620 23624 28626
rect 23572 28562 23624 28568
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23584 27470 23612 28358
rect 23676 27878 23704 29582
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23664 27872 23716 27878
rect 23664 27814 23716 27820
rect 23768 27606 23796 28018
rect 23756 27600 23808 27606
rect 23756 27542 23808 27548
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23584 27010 23612 27406
rect 23584 26982 23704 27010
rect 23570 26888 23626 26897
rect 23204 26852 23256 26858
rect 23570 26823 23572 26832
rect 23204 26794 23256 26800
rect 23624 26823 23626 26832
rect 23572 26794 23624 26800
rect 23112 25424 23164 25430
rect 23112 25366 23164 25372
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 22112 23866 22140 24686
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22112 23322 22140 23598
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 22756 22710 22784 25230
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 21364 22034 21416 22040
rect 21468 22066 21588 22094
rect 21652 22066 21772 22094
rect 21836 22066 21956 22094
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21376 18358 21404 18838
rect 21364 18352 21416 18358
rect 21364 18294 21416 18300
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 14278 21404 14758
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 13734 21404 14214
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21284 12406 21404 12434
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 20904 9454 20956 9460
rect 21008 9438 21128 9466
rect 21180 9512 21232 9518
rect 21232 9472 21312 9500
rect 21180 9454 21232 9460
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20916 9178 20944 9318
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20640 8362 20668 8842
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20732 7478 20760 7754
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20824 7410 20852 7822
rect 21008 7818 21036 9438
rect 21284 9042 21312 9472
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21086 7848 21142 7857
rect 20996 7812 21048 7818
rect 21086 7783 21142 7792
rect 20996 7754 21048 7760
rect 20902 7576 20958 7585
rect 20902 7511 20958 7520
rect 20916 7478 20944 7511
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 6866 20668 7142
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20640 5778 20668 6598
rect 20824 6202 20852 7346
rect 21100 6798 21128 7783
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 20916 6390 20944 6734
rect 21192 6730 21220 8434
rect 21284 6866 21312 8978
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21008 6458 21036 6666
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21100 6202 21128 6258
rect 20824 6174 21128 6202
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20824 5574 20852 6174
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20364 4826 20392 5034
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20732 4049 20760 4082
rect 20718 4040 20774 4049
rect 20076 4004 20128 4010
rect 20718 3975 20774 3984
rect 20076 3946 20128 3952
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3126 14504 3334
rect 16316 3194 16344 3470
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16868 3126 16896 3334
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 18984 3058 19012 3470
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19168 3126 19196 3334
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13556 800 13584 2858
rect 13648 2650 13676 2926
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 14844 800 14872 2926
rect 16684 2650 16712 2926
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16776 800 16804 2858
rect 18064 800 18092 2926
rect 19444 2582 19472 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2450
rect 21192 1714 21220 3538
rect 21376 2774 21404 12406
rect 21468 11778 21496 22066
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21560 18426 21588 18770
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21560 15434 21588 15846
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21560 14822 21588 15370
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21548 14544 21600 14550
rect 21548 14486 21600 14492
rect 21560 13258 21588 14486
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21652 12434 21680 22066
rect 21836 20466 21864 22066
rect 22296 22030 22324 22510
rect 22560 22500 22612 22506
rect 22560 22442 22612 22448
rect 22652 22500 22704 22506
rect 22652 22442 22704 22448
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 22192 20460 22244 20466
rect 22244 20420 22324 20448
rect 22192 20402 22244 20408
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 21744 18698 21772 19110
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 22020 15638 22048 19110
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22112 18358 22140 18702
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 14958 21864 15438
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21732 14884 21784 14890
rect 21732 14826 21784 14832
rect 21744 14618 21772 14826
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21744 13938 21772 14282
rect 21836 14006 21864 14350
rect 21928 14074 21956 14962
rect 22020 14958 22048 15370
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21744 13394 21772 13874
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21836 13394 21864 13738
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21928 13258 21956 14010
rect 22020 13938 22048 14894
rect 22112 14346 22140 16594
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22204 16114 22232 16526
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22204 15502 22232 16050
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22296 15162 22324 20420
rect 22374 19952 22430 19961
rect 22374 19887 22430 19896
rect 22388 19854 22416 19887
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22388 17202 22416 17682
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22376 16720 22428 16726
rect 22376 16662 22428 16668
rect 22388 16538 22416 16662
rect 22480 16658 22508 19382
rect 22572 19174 22600 22442
rect 22664 21486 22692 22442
rect 22756 21962 22784 22646
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22756 21554 22784 21898
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22664 20602 22692 20810
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22572 17338 22600 18294
rect 22664 17678 22692 20402
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22756 18630 22784 20266
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22756 16794 22784 18566
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22388 16510 22508 16538
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22112 13258 22140 14282
rect 22388 13326 22416 16050
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22204 12918 22232 13126
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 21652 12406 21772 12434
rect 21468 11750 21680 11778
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21468 11218 21496 11630
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21560 10849 21588 11086
rect 21546 10840 21602 10849
rect 21546 10775 21602 10784
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21468 8974 21496 9522
rect 21560 9382 21588 10406
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21456 8016 21508 8022
rect 21454 7984 21456 7993
rect 21508 7984 21510 7993
rect 21454 7919 21510 7928
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21468 6798 21496 7414
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21468 6254 21496 6734
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21652 4010 21680 11750
rect 21744 4690 21772 12406
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21928 11898 21956 12174
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22112 10674 22140 11494
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10130 22048 10542
rect 22112 10198 22140 10610
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22020 9110 22048 10066
rect 22112 9518 22140 10134
rect 22204 9994 22232 10950
rect 22296 10810 22324 12786
rect 22388 12434 22416 13262
rect 22480 13190 22508 16510
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22572 14482 22600 15574
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22572 13326 22600 14418
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12594 22508 13126
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22480 12566 22600 12594
rect 22388 12406 22508 12434
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22388 9194 22416 12174
rect 22480 11558 22508 12406
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22480 9586 22508 11290
rect 22572 9654 22600 12566
rect 22664 12434 22692 12786
rect 22664 12406 22784 12434
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 10266 22692 11494
rect 22756 10810 22784 12406
rect 22848 12374 22876 25162
rect 22940 24342 22968 25230
rect 23216 24750 23244 26794
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 23492 25922 23520 26250
rect 23584 26042 23612 26794
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23492 25906 23612 25922
rect 23492 25900 23624 25906
rect 23492 25894 23572 25900
rect 23572 25842 23624 25848
rect 23480 25764 23532 25770
rect 23480 25706 23532 25712
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 22928 24336 22980 24342
rect 22928 24278 22980 24284
rect 22940 18766 22968 24278
rect 23020 24132 23072 24138
rect 23020 24074 23072 24080
rect 23032 22438 23060 24074
rect 23216 22574 23244 24686
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23204 22568 23256 22574
rect 23204 22510 23256 22516
rect 23020 22432 23072 22438
rect 23018 22400 23020 22409
rect 23072 22400 23074 22409
rect 23018 22335 23074 22344
rect 23308 22030 23336 23462
rect 23400 23186 23428 23666
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 23032 19446 23060 21898
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 23124 20058 23152 21490
rect 23296 21412 23348 21418
rect 23296 21354 23348 21360
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23112 20052 23164 20058
rect 23112 19994 23164 20000
rect 23216 19990 23244 20878
rect 23308 20466 23336 21354
rect 23400 20942 23428 22986
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23204 19984 23256 19990
rect 23204 19926 23256 19932
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 23020 19304 23072 19310
rect 23018 19272 23020 19281
rect 23072 19272 23074 19281
rect 23018 19207 23074 19216
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22940 15910 22968 16390
rect 23032 16250 23060 17614
rect 23216 16726 23244 19926
rect 23400 19378 23428 20334
rect 23492 19854 23520 25706
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23584 24410 23612 24686
rect 23572 24404 23624 24410
rect 23572 24346 23624 24352
rect 23676 24206 23704 26982
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 24136 25906 24164 26318
rect 24412 26314 24440 29650
rect 24504 26586 24532 32302
rect 24596 31754 24624 32370
rect 25056 31754 25084 32778
rect 25240 32366 25268 33526
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 24584 31748 24636 31754
rect 24584 31690 24636 31696
rect 25044 31748 25096 31754
rect 25044 31690 25096 31696
rect 24596 31414 24624 31690
rect 25332 31482 25360 36110
rect 25504 35692 25556 35698
rect 25504 35634 25556 35640
rect 25516 34746 25544 35634
rect 25504 34740 25556 34746
rect 25504 34682 25556 34688
rect 25792 34406 25820 36858
rect 25976 36242 26004 37062
rect 25964 36236 26016 36242
rect 25964 36178 26016 36184
rect 26160 35154 26188 37198
rect 26436 36242 26464 39200
rect 27252 37324 27304 37330
rect 27252 37266 27304 37272
rect 26792 36644 26844 36650
rect 26792 36586 26844 36592
rect 26424 36236 26476 36242
rect 26424 36178 26476 36184
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26148 35148 26200 35154
rect 26148 35090 26200 35096
rect 25872 34604 25924 34610
rect 25872 34546 25924 34552
rect 25780 34400 25832 34406
rect 25780 34342 25832 34348
rect 25884 33658 25912 34546
rect 25964 34536 26016 34542
rect 25964 34478 26016 34484
rect 25976 33998 26004 34478
rect 25964 33992 26016 33998
rect 25964 33934 26016 33940
rect 25872 33652 25924 33658
rect 25872 33594 25924 33600
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 25412 33448 25464 33454
rect 25412 33390 25464 33396
rect 25424 31822 25452 33390
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25516 32502 25544 32710
rect 25504 32496 25556 32502
rect 25504 32438 25556 32444
rect 25608 32298 25636 33458
rect 25976 32570 26004 33934
rect 26056 32972 26108 32978
rect 26160 32960 26188 35090
rect 26252 35086 26280 35430
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 26620 34542 26648 34886
rect 26608 34536 26660 34542
rect 26608 34478 26660 34484
rect 26240 33992 26292 33998
rect 26240 33934 26292 33940
rect 26252 33658 26280 33934
rect 26700 33924 26752 33930
rect 26700 33866 26752 33872
rect 26332 33856 26384 33862
rect 26332 33798 26384 33804
rect 26240 33652 26292 33658
rect 26240 33594 26292 33600
rect 26344 32978 26372 33798
rect 26108 32932 26188 32960
rect 26056 32914 26108 32920
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 25872 32496 25924 32502
rect 25872 32438 25924 32444
rect 25688 32360 25740 32366
rect 25688 32302 25740 32308
rect 25596 32292 25648 32298
rect 25596 32234 25648 32240
rect 25412 31816 25464 31822
rect 25412 31758 25464 31764
rect 25320 31476 25372 31482
rect 25320 31418 25372 31424
rect 25424 31414 25452 31758
rect 25700 31754 25728 32302
rect 25700 31726 25820 31754
rect 24584 31408 24636 31414
rect 24584 31350 24636 31356
rect 25412 31408 25464 31414
rect 25412 31350 25464 31356
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 24952 30660 25004 30666
rect 24952 30602 25004 30608
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24872 29850 24900 30194
rect 24964 30190 24992 30602
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24780 29306 24808 29446
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 25056 29238 25084 31282
rect 25136 30728 25188 30734
rect 25136 30670 25188 30676
rect 24676 29232 24728 29238
rect 24676 29174 24728 29180
rect 25044 29232 25096 29238
rect 25044 29174 25096 29180
rect 24688 27470 24716 29174
rect 25148 29034 25176 30670
rect 25320 30592 25372 30598
rect 25320 30534 25372 30540
rect 25136 29028 25188 29034
rect 25136 28970 25188 28976
rect 25148 28762 25176 28970
rect 25136 28756 25188 28762
rect 25136 28698 25188 28704
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 24768 27872 24820 27878
rect 24768 27814 24820 27820
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24492 26580 24544 26586
rect 24492 26522 24544 26528
rect 24400 26308 24452 26314
rect 24400 26250 24452 26256
rect 24596 25906 24624 27338
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24688 27062 24716 27270
rect 24676 27056 24728 27062
rect 24676 26998 24728 27004
rect 24780 26382 24808 27814
rect 24860 27056 24912 27062
rect 24860 26998 24912 27004
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24872 26042 24900 26998
rect 25148 26926 25176 27950
rect 25332 27946 25360 30534
rect 25424 29850 25452 31350
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 25424 29646 25452 29786
rect 25412 29640 25464 29646
rect 25412 29582 25464 29588
rect 25502 29336 25558 29345
rect 25502 29271 25558 29280
rect 25516 29238 25544 29271
rect 25504 29232 25556 29238
rect 25504 29174 25556 29180
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25320 27940 25372 27946
rect 25320 27882 25372 27888
rect 25136 26920 25188 26926
rect 25136 26862 25188 26868
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 24124 25900 24176 25906
rect 24124 25842 24176 25848
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 24032 24880 24084 24886
rect 24032 24822 24084 24828
rect 24044 24342 24072 24822
rect 24032 24336 24084 24342
rect 24032 24278 24084 24284
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23676 23662 23704 24142
rect 24136 23866 24164 25842
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23768 23526 23796 23802
rect 24688 23730 24716 23802
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23584 22166 23612 22510
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23572 22160 23624 22166
rect 23572 22102 23624 22108
rect 23584 21010 23612 22102
rect 23676 22030 23704 22442
rect 23860 22094 23888 23666
rect 24596 23254 24624 23666
rect 24584 23248 24636 23254
rect 24584 23190 24636 23196
rect 24596 23050 24624 23190
rect 24584 23044 24636 23050
rect 24584 22986 24636 22992
rect 24308 22976 24360 22982
rect 24308 22918 24360 22924
rect 24492 22976 24544 22982
rect 24688 22930 24716 23666
rect 24544 22924 24716 22930
rect 24492 22918 24716 22924
rect 24320 22778 24348 22918
rect 24504 22902 24716 22918
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 23768 22066 23888 22094
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23768 21842 23796 22066
rect 23938 21992 23994 22001
rect 23938 21927 23994 21936
rect 23848 21888 23900 21894
rect 23768 21836 23848 21842
rect 23768 21830 23900 21836
rect 23768 21814 23888 21830
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23572 20868 23624 20874
rect 23572 20810 23624 20816
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23308 18766 23336 19110
rect 23400 18902 23428 19314
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23492 17882 23520 19790
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23204 16584 23256 16590
rect 23202 16552 23204 16561
rect 23256 16552 23258 16561
rect 23112 16516 23164 16522
rect 23202 16487 23258 16496
rect 23112 16458 23164 16464
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23124 16114 23152 16458
rect 23308 16454 23336 17614
rect 23584 17610 23612 20810
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 20534 23704 20742
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23768 20398 23796 21286
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23860 20262 23888 20946
rect 23952 20942 23980 21927
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24412 21622 24440 21830
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22940 12918 22968 15846
rect 23216 15638 23244 16118
rect 23204 15632 23256 15638
rect 23204 15574 23256 15580
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23308 14618 23336 14962
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23584 14482 23612 15098
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23308 13870 23336 14418
rect 23676 14346 23704 18906
rect 23768 17882 23796 19246
rect 23860 18358 23888 19654
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23860 17678 23888 18022
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23860 17270 23888 17478
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23216 13530 23244 13806
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23400 13326 23428 14214
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23020 13252 23072 13258
rect 23020 13194 23072 13200
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 22940 12238 22968 12718
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 22940 11150 22968 11290
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 22756 10554 22784 10746
rect 22756 10526 22876 10554
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22756 10130 22784 10406
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22112 9178 22416 9194
rect 22100 9172 22416 9178
rect 22152 9166 22416 9172
rect 22100 9114 22152 9120
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 22192 8968 22244 8974
rect 22284 8968 22336 8974
rect 22192 8910 22244 8916
rect 22282 8936 22284 8945
rect 22336 8936 22338 8945
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22020 7410 22048 8434
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22020 6798 22048 7346
rect 22112 7342 22140 7958
rect 22204 7954 22232 8910
rect 22282 8871 22338 8880
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22204 7546 22232 7890
rect 22388 7886 22416 8230
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22388 7478 22416 7822
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22112 6780 22140 7278
rect 22192 6792 22244 6798
rect 22112 6752 22192 6780
rect 22020 5914 22048 6734
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 22112 4826 22140 6752
rect 22192 6734 22244 6740
rect 22480 6662 22508 8842
rect 22664 8090 22692 9862
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22756 9178 22784 9318
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22848 9058 22876 10526
rect 22940 9110 22968 11086
rect 22756 9030 22876 9058
rect 22928 9104 22980 9110
rect 22928 9046 22980 9052
rect 22756 8838 22784 9030
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22848 8634 22876 8910
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22836 8492 22888 8498
rect 22888 8452 22968 8480
rect 22836 8434 22888 8440
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22940 7818 22968 8452
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 23032 7562 23060 13194
rect 23308 12866 23336 13194
rect 23308 12850 23428 12866
rect 23308 12844 23440 12850
rect 23308 12838 23388 12844
rect 23388 12786 23440 12792
rect 23492 12646 23520 13194
rect 23952 12918 23980 20878
rect 24504 19854 24532 21286
rect 24596 21010 24624 21830
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24136 16130 24164 19722
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24228 18290 24256 18906
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18358 24624 18566
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24596 16998 24624 17478
rect 24688 17338 24716 22902
rect 24780 21622 24808 25230
rect 25424 24750 25452 25638
rect 25516 25498 25544 25842
rect 25608 25770 25636 29106
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25700 26790 25728 27406
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25596 25764 25648 25770
rect 25596 25706 25648 25712
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25608 25294 25636 25706
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25148 24206 25176 24550
rect 25424 24206 25452 24686
rect 25792 24274 25820 31726
rect 25884 31686 25912 32438
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26068 31822 26096 32370
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 25872 31680 25924 31686
rect 25872 31622 25924 31628
rect 26068 31346 26096 31758
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 26160 31210 26188 32932
rect 26332 32972 26384 32978
rect 26332 32914 26384 32920
rect 26424 32972 26476 32978
rect 26424 32914 26476 32920
rect 26436 32774 26464 32914
rect 26424 32768 26476 32774
rect 26424 32710 26476 32716
rect 26424 32496 26476 32502
rect 26424 32438 26476 32444
rect 25872 31204 25924 31210
rect 25872 31146 25924 31152
rect 26148 31204 26200 31210
rect 26148 31146 26200 31152
rect 25884 30938 25912 31146
rect 25872 30932 25924 30938
rect 25872 30874 25924 30880
rect 26160 30802 26188 31146
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 26160 30138 26188 30738
rect 26240 30184 26292 30190
rect 26160 30132 26240 30138
rect 26160 30126 26292 30132
rect 26160 30110 26280 30126
rect 26436 30122 26464 32438
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26608 31340 26660 31346
rect 26608 31282 26660 31288
rect 26424 30116 26476 30122
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 26068 29170 26096 29514
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 26068 29073 26096 29106
rect 26054 29064 26110 29073
rect 25964 29028 26016 29034
rect 26054 28999 26110 29008
rect 25964 28970 26016 28976
rect 25872 28484 25924 28490
rect 25872 28426 25924 28432
rect 25884 28218 25912 28426
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 25884 25226 25912 26522
rect 25976 26450 26004 28970
rect 26160 28626 26188 30110
rect 26424 30058 26476 30064
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 26068 27470 26096 28018
rect 26252 28014 26280 28902
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 26344 28082 26372 28358
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 26436 27860 26464 30058
rect 26528 29102 26556 31282
rect 26620 30054 26648 31282
rect 26608 30048 26660 30054
rect 26608 29990 26660 29996
rect 26620 29578 26648 29990
rect 26608 29572 26660 29578
rect 26608 29514 26660 29520
rect 26712 29510 26740 33866
rect 26804 31754 26832 36586
rect 27264 35834 27292 37266
rect 28264 36780 28316 36786
rect 28264 36722 28316 36728
rect 27804 36576 27856 36582
rect 27804 36518 27856 36524
rect 27988 36576 28040 36582
rect 27988 36518 28040 36524
rect 27252 35828 27304 35834
rect 27252 35770 27304 35776
rect 27816 35698 27844 36518
rect 26976 35692 27028 35698
rect 26976 35634 27028 35640
rect 27344 35692 27396 35698
rect 27344 35634 27396 35640
rect 27804 35692 27856 35698
rect 27804 35634 27856 35640
rect 26884 35488 26936 35494
rect 26884 35430 26936 35436
rect 26896 34678 26924 35430
rect 26884 34672 26936 34678
rect 26884 34614 26936 34620
rect 26988 34134 27016 35634
rect 27356 35290 27384 35634
rect 28000 35630 28028 36518
rect 27988 35624 28040 35630
rect 27988 35566 28040 35572
rect 28276 35442 28304 36722
rect 28368 35630 28396 39200
rect 29656 38026 29684 39200
rect 29656 37998 29776 38026
rect 29552 37188 29604 37194
rect 29552 37130 29604 37136
rect 29644 37188 29696 37194
rect 29644 37130 29696 37136
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28540 36168 28592 36174
rect 28540 36110 28592 36116
rect 28448 36032 28500 36038
rect 28448 35974 28500 35980
rect 28356 35624 28408 35630
rect 28356 35566 28408 35572
rect 28276 35414 28396 35442
rect 27344 35284 27396 35290
rect 27344 35226 27396 35232
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 28264 35080 28316 35086
rect 28264 35022 28316 35028
rect 27344 34400 27396 34406
rect 27344 34342 27396 34348
rect 26976 34128 27028 34134
rect 26976 34070 27028 34076
rect 26988 33522 27016 34070
rect 27356 34066 27384 34342
rect 27344 34060 27396 34066
rect 27344 34002 27396 34008
rect 27540 33862 27568 35022
rect 27712 34672 27764 34678
rect 27712 34614 27764 34620
rect 27724 33998 27752 34614
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 26988 32570 27016 33458
rect 27068 33312 27120 33318
rect 27068 33254 27120 33260
rect 27080 32842 27108 33254
rect 27068 32836 27120 32842
rect 27068 32778 27120 32784
rect 26976 32564 27028 32570
rect 26976 32506 27028 32512
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 26804 31726 26924 31754
rect 26792 31680 26844 31686
rect 26792 31622 26844 31628
rect 26804 30598 26832 31622
rect 26792 30592 26844 30598
rect 26792 30534 26844 30540
rect 26804 29850 26832 30534
rect 26792 29844 26844 29850
rect 26792 29786 26844 29792
rect 26896 29594 26924 31726
rect 27080 31414 27108 32370
rect 27724 32298 27752 33934
rect 27896 33924 27948 33930
rect 27896 33866 27948 33872
rect 27908 33522 27936 33866
rect 28184 33522 28212 34546
rect 28276 34474 28304 35022
rect 28264 34468 28316 34474
rect 28264 34410 28316 34416
rect 27896 33516 27948 33522
rect 27896 33458 27948 33464
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27988 33448 28040 33454
rect 27988 33390 28040 33396
rect 27816 32570 27844 33390
rect 27896 32972 27948 32978
rect 27896 32914 27948 32920
rect 27804 32564 27856 32570
rect 27804 32506 27856 32512
rect 27712 32292 27764 32298
rect 27712 32234 27764 32240
rect 27344 32224 27396 32230
rect 27344 32166 27396 32172
rect 27068 31408 27120 31414
rect 27068 31350 27120 31356
rect 27080 30598 27108 31350
rect 27160 31136 27212 31142
rect 27160 31078 27212 31084
rect 27068 30592 27120 30598
rect 27068 30534 27120 30540
rect 26974 29880 27030 29889
rect 26974 29815 26976 29824
rect 27028 29815 27030 29824
rect 26976 29786 27028 29792
rect 26804 29566 26924 29594
rect 26700 29504 26752 29510
rect 26700 29446 26752 29452
rect 26516 29096 26568 29102
rect 26516 29038 26568 29044
rect 26804 27860 26832 29566
rect 26988 29170 27016 29786
rect 27080 29322 27108 30534
rect 27172 30394 27200 31078
rect 27160 30388 27212 30394
rect 27160 30330 27212 30336
rect 27252 30320 27304 30326
rect 27250 30288 27252 30297
rect 27304 30288 27306 30297
rect 27250 30223 27306 30232
rect 27252 30048 27304 30054
rect 27252 29990 27304 29996
rect 27080 29306 27200 29322
rect 27080 29300 27212 29306
rect 27080 29294 27160 29300
rect 27160 29242 27212 29248
rect 27264 29238 27292 29990
rect 27356 29646 27384 32166
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27436 30320 27488 30326
rect 27436 30262 27488 30268
rect 27448 30054 27476 30262
rect 27540 30054 27568 31826
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27528 30048 27580 30054
rect 27528 29990 27580 29996
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27540 29578 27568 29990
rect 27632 29646 27660 31758
rect 27804 31748 27856 31754
rect 27804 31690 27856 31696
rect 27816 31482 27844 31690
rect 27804 31476 27856 31482
rect 27804 31418 27856 31424
rect 27712 30320 27764 30326
rect 27710 30288 27712 30297
rect 27764 30288 27766 30297
rect 27710 30223 27766 30232
rect 27908 30122 27936 32914
rect 28000 32230 28028 33390
rect 28184 33114 28212 33458
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 28184 32502 28212 33050
rect 28172 32496 28224 32502
rect 28172 32438 28224 32444
rect 27988 32224 28040 32230
rect 27988 32166 28040 32172
rect 28368 32178 28396 35414
rect 28460 35018 28488 35974
rect 28552 35290 28580 36110
rect 28540 35284 28592 35290
rect 28540 35226 28592 35232
rect 28552 35086 28580 35226
rect 28540 35080 28592 35086
rect 28540 35022 28592 35028
rect 28448 35012 28500 35018
rect 28448 34954 28500 34960
rect 28552 34678 28580 35022
rect 28632 34740 28684 34746
rect 28632 34682 28684 34688
rect 28540 34672 28592 34678
rect 28540 34614 28592 34620
rect 28540 34536 28592 34542
rect 28540 34478 28592 34484
rect 28552 33114 28580 34478
rect 28540 33108 28592 33114
rect 28540 33050 28592 33056
rect 28552 32910 28580 33050
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28448 32768 28500 32774
rect 28448 32710 28500 32716
rect 28460 32298 28488 32710
rect 28448 32292 28500 32298
rect 28448 32234 28500 32240
rect 28644 32230 28672 34682
rect 28736 34610 28764 37062
rect 29000 36712 29052 36718
rect 29000 36654 29052 36660
rect 29012 36174 29040 36654
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 28816 36100 28868 36106
rect 28816 36042 28868 36048
rect 28828 34610 28856 36042
rect 29564 35834 29592 37130
rect 29656 36378 29684 37130
rect 29748 36650 29776 37998
rect 30944 37194 30972 39200
rect 30932 37188 30984 37194
rect 30932 37130 30984 37136
rect 30196 36712 30248 36718
rect 30196 36654 30248 36660
rect 29736 36644 29788 36650
rect 29736 36586 29788 36592
rect 30208 36378 30236 36654
rect 31668 36576 31720 36582
rect 31668 36518 31720 36524
rect 29644 36372 29696 36378
rect 29644 36314 29696 36320
rect 30196 36372 30248 36378
rect 30196 36314 30248 36320
rect 31680 36242 31708 36518
rect 32232 36242 32260 39200
rect 32876 36718 32904 39200
rect 36740 37618 36768 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 36740 37590 36860 37618
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 36726 37496 36782 37505
rect 36726 37431 36782 37440
rect 34888 37392 34940 37398
rect 34888 37334 34940 37340
rect 34796 37188 34848 37194
rect 34796 37130 34848 37136
rect 32404 36712 32456 36718
rect 32404 36654 32456 36660
rect 32588 36712 32640 36718
rect 32588 36654 32640 36660
rect 32864 36712 32916 36718
rect 32864 36654 32916 36660
rect 31668 36236 31720 36242
rect 31668 36178 31720 36184
rect 32220 36236 32272 36242
rect 32220 36178 32272 36184
rect 31852 36100 31904 36106
rect 31852 36042 31904 36048
rect 31864 35834 31892 36042
rect 29552 35828 29604 35834
rect 29552 35770 29604 35776
rect 31852 35828 31904 35834
rect 31852 35770 31904 35776
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 32220 35692 32272 35698
rect 32220 35634 32272 35640
rect 29000 35080 29052 35086
rect 29000 35022 29052 35028
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29012 34746 29040 35022
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 28724 34604 28776 34610
rect 28724 34546 28776 34552
rect 28816 34604 28868 34610
rect 28816 34546 28868 34552
rect 28736 34066 28764 34546
rect 29000 34536 29052 34542
rect 29000 34478 29052 34484
rect 29012 34202 29040 34478
rect 29932 34202 29960 35022
rect 29000 34196 29052 34202
rect 29000 34138 29052 34144
rect 29920 34196 29972 34202
rect 29920 34138 29972 34144
rect 30116 34134 30144 35634
rect 31300 35080 31352 35086
rect 31300 35022 31352 35028
rect 31116 34740 31168 34746
rect 31312 34728 31340 35022
rect 31392 34944 31444 34950
rect 31392 34886 31444 34892
rect 31404 34746 31432 34886
rect 31168 34700 31340 34728
rect 31116 34682 31168 34688
rect 30656 34400 30708 34406
rect 30656 34342 30708 34348
rect 30748 34400 30800 34406
rect 30748 34342 30800 34348
rect 30104 34128 30156 34134
rect 30104 34070 30156 34076
rect 28724 34060 28776 34066
rect 28724 34002 28776 34008
rect 29920 33992 29972 33998
rect 29920 33934 29972 33940
rect 30564 33992 30616 33998
rect 30564 33934 30616 33940
rect 29000 33312 29052 33318
rect 29000 33254 29052 33260
rect 29012 32910 29040 33254
rect 28724 32904 28776 32910
rect 28724 32846 28776 32852
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 29828 32904 29880 32910
rect 29828 32846 29880 32852
rect 28632 32224 28684 32230
rect 28000 31890 28028 32166
rect 28368 32150 28580 32178
rect 28632 32166 28684 32172
rect 28172 31952 28224 31958
rect 28172 31894 28224 31900
rect 27988 31884 28040 31890
rect 27988 31826 28040 31832
rect 27988 30660 28040 30666
rect 27988 30602 28040 30608
rect 27896 30116 27948 30122
rect 27896 30058 27948 30064
rect 27712 29776 27764 29782
rect 27712 29718 27764 29724
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27528 29572 27580 29578
rect 27528 29514 27580 29520
rect 27724 29306 27752 29718
rect 27908 29578 27936 30058
rect 28000 29850 28028 30602
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 28092 29889 28120 30194
rect 28078 29880 28134 29889
rect 27988 29844 28040 29850
rect 28078 29815 28134 29824
rect 27988 29786 28040 29792
rect 28184 29782 28212 31894
rect 28552 31754 28580 32150
rect 28552 31726 28672 31754
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 28368 31346 28396 31622
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28368 30802 28396 31282
rect 28540 31136 28592 31142
rect 28540 31078 28592 31084
rect 28356 30796 28408 30802
rect 28356 30738 28408 30744
rect 28264 30592 28316 30598
rect 28264 30534 28316 30540
rect 28276 29850 28304 30534
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28172 29776 28224 29782
rect 28172 29718 28224 29724
rect 27896 29572 27948 29578
rect 27896 29514 27948 29520
rect 27712 29300 27764 29306
rect 27712 29242 27764 29248
rect 27252 29232 27304 29238
rect 27252 29174 27304 29180
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 27160 29164 27212 29170
rect 27160 29106 27212 29112
rect 26988 28994 27016 29106
rect 26896 28966 27016 28994
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 26896 28694 26924 28966
rect 26884 28688 26936 28694
rect 26884 28630 26936 28636
rect 26884 28552 26936 28558
rect 26884 28494 26936 28500
rect 26896 27946 26924 28494
rect 26884 27940 26936 27946
rect 26884 27882 26936 27888
rect 26252 27832 26464 27860
rect 26712 27832 26832 27860
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 26056 26376 26108 26382
rect 26108 26336 26188 26364
rect 26056 26318 26108 26324
rect 25964 26240 26016 26246
rect 25964 26182 26016 26188
rect 25976 25838 26004 26182
rect 26160 25838 26188 26336
rect 25964 25832 26016 25838
rect 25964 25774 26016 25780
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 25872 25220 25924 25226
rect 25872 25162 25924 25168
rect 26160 24750 26188 25774
rect 26148 24744 26200 24750
rect 26068 24692 26148 24698
rect 26068 24686 26200 24692
rect 25964 24676 26016 24682
rect 26068 24670 26188 24686
rect 26068 24664 26096 24670
rect 26016 24636 26096 24664
rect 25964 24618 26016 24624
rect 26148 24608 26200 24614
rect 26148 24550 26200 24556
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25608 23254 25636 23598
rect 25596 23248 25648 23254
rect 25596 23190 25648 23196
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24964 21962 24992 22986
rect 25056 22234 25084 23054
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 24768 21616 24820 21622
rect 24768 21558 24820 21564
rect 25424 21418 25452 23054
rect 25792 23050 25820 24210
rect 26160 24206 26188 24550
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 25780 23044 25832 23050
rect 25780 22986 25832 22992
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25516 22710 25544 22918
rect 25504 22704 25556 22710
rect 25504 22646 25556 22652
rect 26160 22506 26188 24142
rect 26252 23186 26280 27832
rect 26332 27464 26384 27470
rect 26330 27432 26332 27441
rect 26384 27432 26386 27441
rect 26330 27367 26386 27376
rect 26424 26376 26476 26382
rect 26424 26318 26476 26324
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26344 25906 26372 26250
rect 26436 25974 26464 26318
rect 26424 25968 26476 25974
rect 26424 25910 26476 25916
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26332 25152 26384 25158
rect 26332 25094 26384 25100
rect 26344 24138 26372 25094
rect 26712 24682 26740 27832
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26804 26586 26832 27406
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 26896 25158 26924 27882
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 26988 25702 27016 27406
rect 27080 25974 27108 28970
rect 27172 28490 27200 29106
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27252 28960 27304 28966
rect 27252 28902 27304 28908
rect 27264 28558 27292 28902
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27160 28484 27212 28490
rect 27160 28426 27212 28432
rect 27172 28082 27200 28426
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27436 28144 27488 28150
rect 27436 28086 27488 28092
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27344 27600 27396 27606
rect 27342 27568 27344 27577
rect 27396 27568 27398 27577
rect 27342 27503 27398 27512
rect 27448 27402 27476 28086
rect 27540 28082 27568 28358
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27528 27600 27580 27606
rect 27528 27542 27580 27548
rect 27540 27470 27568 27542
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27436 27396 27488 27402
rect 27436 27338 27488 27344
rect 27448 27305 27476 27338
rect 27434 27296 27490 27305
rect 27434 27231 27490 27240
rect 27540 27130 27568 27406
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 27540 26314 27568 27066
rect 27528 26308 27580 26314
rect 27528 26250 27580 26256
rect 27068 25968 27120 25974
rect 27068 25910 27120 25916
rect 26976 25696 27028 25702
rect 26976 25638 27028 25644
rect 27080 25294 27108 25910
rect 27252 25492 27304 25498
rect 27252 25434 27304 25440
rect 27068 25288 27120 25294
rect 27068 25230 27120 25236
rect 26884 25152 26936 25158
rect 26884 25094 26936 25100
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 26700 24676 26752 24682
rect 26700 24618 26752 24624
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26436 24274 26464 24550
rect 27172 24410 27200 24754
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 26332 24132 26384 24138
rect 26332 24074 26384 24080
rect 27264 23866 27292 25434
rect 27632 25294 27660 29038
rect 27908 28150 27936 29514
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 27896 28144 27948 28150
rect 27896 28086 27948 28092
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27804 27464 27856 27470
rect 27804 27406 27856 27412
rect 27894 27432 27950 27441
rect 27724 26926 27752 27406
rect 27712 26920 27764 26926
rect 27712 26862 27764 26868
rect 27816 26518 27844 27406
rect 27894 27367 27950 27376
rect 27908 27334 27936 27367
rect 27896 27328 27948 27334
rect 27896 27270 27948 27276
rect 27804 26512 27856 26518
rect 27804 26454 27856 26460
rect 28000 26382 28028 29446
rect 28446 29336 28502 29345
rect 28446 29271 28448 29280
rect 28500 29271 28502 29280
rect 28448 29242 28500 29248
rect 28552 29170 28580 31078
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 28184 27674 28488 27690
rect 28172 27668 28500 27674
rect 28224 27662 28448 27668
rect 28172 27610 28224 27616
rect 28448 27610 28500 27616
rect 28170 27568 28226 27577
rect 28080 27532 28132 27538
rect 28170 27503 28172 27512
rect 28080 27474 28132 27480
rect 28224 27503 28226 27512
rect 28172 27474 28224 27480
rect 27988 26376 28040 26382
rect 27988 26318 28040 26324
rect 27896 26308 27948 26314
rect 27896 26250 27948 26256
rect 27908 26042 27936 26250
rect 27896 26036 27948 26042
rect 27896 25978 27948 25984
rect 28092 25770 28120 27474
rect 28448 27464 28500 27470
rect 28448 27406 28500 27412
rect 28354 27296 28410 27305
rect 28354 27231 28410 27240
rect 28368 26858 28396 27231
rect 28356 26852 28408 26858
rect 28356 26794 28408 26800
rect 28460 26790 28488 27406
rect 28448 26784 28500 26790
rect 28448 26726 28500 26732
rect 28460 26450 28488 26726
rect 28540 26512 28592 26518
rect 28540 26454 28592 26460
rect 28448 26444 28500 26450
rect 28448 26386 28500 26392
rect 28080 25764 28132 25770
rect 28080 25706 28132 25712
rect 27896 25696 27948 25702
rect 27896 25638 27948 25644
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27908 25226 27936 25638
rect 27896 25220 27948 25226
rect 27896 25162 27948 25168
rect 27344 25152 27396 25158
rect 27804 25152 27856 25158
rect 27344 25094 27396 25100
rect 27724 25112 27804 25140
rect 27356 24954 27384 25094
rect 27344 24948 27396 24954
rect 27344 24890 27396 24896
rect 27724 24750 27752 25112
rect 27804 25094 27856 25100
rect 27712 24744 27764 24750
rect 27712 24686 27764 24692
rect 27908 24410 27936 25162
rect 28448 24880 28500 24886
rect 28448 24822 28500 24828
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 28368 24410 28396 24686
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 28356 24404 28408 24410
rect 28356 24346 28408 24352
rect 27436 24132 27488 24138
rect 27436 24074 27488 24080
rect 27448 23866 27476 24074
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27436 23860 27488 23866
rect 27436 23802 27488 23808
rect 26332 23792 26384 23798
rect 26332 23734 26384 23740
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26148 22500 26200 22506
rect 26148 22442 26200 22448
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 25516 22030 25544 22374
rect 26160 22098 26188 22442
rect 26148 22092 26200 22098
rect 26344 22094 26372 23734
rect 28460 23225 28488 24822
rect 28552 24206 28580 26454
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28644 24154 28672 31726
rect 28736 31278 28764 32846
rect 28908 32564 28960 32570
rect 28908 32506 28960 32512
rect 28816 32224 28868 32230
rect 28816 32166 28868 32172
rect 28724 31272 28776 31278
rect 28724 31214 28776 31220
rect 28828 29578 28856 32166
rect 28920 30666 28948 32506
rect 29840 32502 29868 32846
rect 29184 32496 29236 32502
rect 29736 32496 29788 32502
rect 29184 32438 29236 32444
rect 29734 32464 29736 32473
rect 29828 32496 29880 32502
rect 29788 32464 29790 32473
rect 29092 32020 29144 32026
rect 29092 31962 29144 31968
rect 29104 31754 29132 31962
rect 29196 31958 29224 32438
rect 29828 32438 29880 32444
rect 29734 32399 29790 32408
rect 29184 31952 29236 31958
rect 29184 31894 29236 31900
rect 29012 31726 29132 31754
rect 28908 30660 28960 30666
rect 28908 30602 28960 30608
rect 29012 30326 29040 31726
rect 29196 31142 29224 31894
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 29184 31136 29236 31142
rect 29184 31078 29236 31084
rect 29196 30734 29224 31078
rect 29184 30728 29236 30734
rect 29184 30670 29236 30676
rect 29840 30666 29868 31826
rect 29932 31822 29960 33934
rect 30012 33856 30064 33862
rect 30012 33798 30064 33804
rect 30024 33590 30052 33798
rect 30012 33584 30064 33590
rect 30012 33526 30064 33532
rect 30196 33584 30248 33590
rect 30196 33526 30248 33532
rect 30208 33114 30236 33526
rect 30196 33108 30248 33114
rect 30196 33050 30248 33056
rect 30472 32972 30524 32978
rect 30472 32914 30524 32920
rect 30104 32904 30156 32910
rect 30484 32881 30512 32914
rect 30104 32846 30156 32852
rect 30470 32872 30526 32881
rect 30116 32570 30144 32846
rect 30470 32807 30526 32816
rect 30104 32564 30156 32570
rect 30104 32506 30156 32512
rect 30196 32428 30248 32434
rect 30196 32370 30248 32376
rect 30288 32428 30340 32434
rect 30288 32370 30340 32376
rect 29920 31816 29972 31822
rect 29920 31758 29972 31764
rect 30208 31754 30236 32370
rect 30300 32026 30328 32370
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 30116 31726 30236 31754
rect 29920 31680 29972 31686
rect 29920 31622 29972 31628
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 29932 31414 29960 31622
rect 29920 31408 29972 31414
rect 29920 31350 29972 31356
rect 29920 31136 29972 31142
rect 29920 31078 29972 31084
rect 29932 30734 29960 31078
rect 29920 30728 29972 30734
rect 29920 30670 29972 30676
rect 29828 30660 29880 30666
rect 29828 30602 29880 30608
rect 29184 30388 29236 30394
rect 29184 30330 29236 30336
rect 29000 30320 29052 30326
rect 29052 30268 29132 30274
rect 29000 30262 29132 30268
rect 29012 30246 29132 30262
rect 29000 30116 29052 30122
rect 29000 30058 29052 30064
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 28816 29572 28868 29578
rect 28816 29514 28868 29520
rect 28828 29322 28856 29514
rect 28736 29294 28856 29322
rect 28736 29034 28764 29294
rect 28816 29164 28868 29170
rect 28816 29106 28868 29112
rect 28724 29028 28776 29034
rect 28724 28970 28776 28976
rect 28736 28762 28764 28970
rect 28724 28756 28776 28762
rect 28724 28698 28776 28704
rect 28724 27940 28776 27946
rect 28724 27882 28776 27888
rect 28736 26450 28764 27882
rect 28828 27606 28856 29106
rect 28920 29034 28948 29786
rect 28908 29028 28960 29034
rect 28908 28970 28960 28976
rect 29012 28762 29040 30058
rect 29104 29510 29132 30246
rect 29092 29504 29144 29510
rect 29092 29446 29144 29452
rect 29196 29238 29224 30330
rect 29276 30116 29328 30122
rect 29276 30058 29328 30064
rect 29288 29850 29316 30058
rect 29276 29844 29328 29850
rect 29276 29786 29328 29792
rect 29184 29232 29236 29238
rect 29184 29174 29236 29180
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29840 28694 29868 30602
rect 30024 30394 30052 31622
rect 30012 30388 30064 30394
rect 30012 30330 30064 30336
rect 30116 30274 30144 31726
rect 30300 31464 30328 31826
rect 30576 31754 30604 33934
rect 30668 33114 30696 34342
rect 30760 33114 30788 34342
rect 31312 33998 31340 34700
rect 31392 34740 31444 34746
rect 31392 34682 31444 34688
rect 30932 33992 30984 33998
rect 30932 33934 30984 33940
rect 31300 33992 31352 33998
rect 31300 33934 31352 33940
rect 30944 33454 30972 33934
rect 32128 33856 32180 33862
rect 32128 33798 32180 33804
rect 32140 33522 32168 33798
rect 32128 33516 32180 33522
rect 32128 33458 32180 33464
rect 30932 33448 30984 33454
rect 30932 33390 30984 33396
rect 31024 33448 31076 33454
rect 31024 33390 31076 33396
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30748 33108 30800 33114
rect 30748 33050 30800 33056
rect 30760 32994 30788 33050
rect 30668 32966 30788 32994
rect 30668 32570 30696 32966
rect 30852 32910 30880 33254
rect 30840 32904 30892 32910
rect 30840 32846 30892 32852
rect 30656 32564 30708 32570
rect 30656 32506 30708 32512
rect 30472 31748 30604 31754
rect 30524 31726 30604 31748
rect 30472 31690 30524 31696
rect 30380 31476 30432 31482
rect 30300 31436 30380 31464
rect 30380 31418 30432 31424
rect 30668 31414 30696 32506
rect 30748 32292 30800 32298
rect 30748 32234 30800 32240
rect 30760 32065 30788 32234
rect 30746 32056 30802 32065
rect 30746 31991 30802 32000
rect 30840 31884 30892 31890
rect 30840 31826 30892 31832
rect 30656 31408 30708 31414
rect 30656 31350 30708 31356
rect 30656 31272 30708 31278
rect 30656 31214 30708 31220
rect 30668 30938 30696 31214
rect 30656 30932 30708 30938
rect 30656 30874 30708 30880
rect 30196 30728 30248 30734
rect 30196 30670 30248 30676
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30024 30246 30144 30274
rect 29920 29776 29972 29782
rect 29920 29718 29972 29724
rect 29932 29306 29960 29718
rect 29920 29300 29972 29306
rect 29920 29242 29972 29248
rect 29828 28688 29880 28694
rect 29828 28630 29880 28636
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29012 28098 29040 28358
rect 29840 28150 29868 28494
rect 28920 28082 29040 28098
rect 29828 28144 29880 28150
rect 29828 28086 29880 28092
rect 28920 28076 29052 28082
rect 28920 28070 29000 28076
rect 28816 27600 28868 27606
rect 28816 27542 28868 27548
rect 28920 27418 28948 28070
rect 29000 28018 29052 28024
rect 30024 28014 30052 30246
rect 30104 30184 30156 30190
rect 30104 30126 30156 30132
rect 30116 29850 30144 30126
rect 30104 29844 30156 29850
rect 30104 29786 30156 29792
rect 30208 28422 30236 30670
rect 30288 30660 30340 30666
rect 30288 30602 30340 30608
rect 30300 30394 30328 30602
rect 30288 30388 30340 30394
rect 30288 30330 30340 30336
rect 30300 29782 30328 30330
rect 30392 30326 30420 30670
rect 30748 30660 30800 30666
rect 30748 30602 30800 30608
rect 30472 30592 30524 30598
rect 30472 30534 30524 30540
rect 30380 30320 30432 30326
rect 30380 30262 30432 30268
rect 30288 29776 30340 29782
rect 30288 29718 30340 29724
rect 30484 29084 30512 30534
rect 30760 30433 30788 30602
rect 30746 30424 30802 30433
rect 30746 30359 30802 30368
rect 30852 30326 30880 31826
rect 30944 31278 30972 33390
rect 31036 33046 31064 33390
rect 31760 33312 31812 33318
rect 31760 33254 31812 33260
rect 32036 33312 32088 33318
rect 32036 33254 32088 33260
rect 31772 33114 31800 33254
rect 31576 33108 31628 33114
rect 31576 33050 31628 33056
rect 31760 33108 31812 33114
rect 31760 33050 31812 33056
rect 31852 33108 31904 33114
rect 31852 33050 31904 33056
rect 31024 33040 31076 33046
rect 31024 32982 31076 32988
rect 31300 32904 31352 32910
rect 31024 32882 31076 32888
rect 31024 32824 31076 32830
rect 31298 32872 31300 32881
rect 31352 32872 31354 32881
rect 31036 31396 31064 32824
rect 31588 32842 31616 33050
rect 31298 32807 31354 32816
rect 31576 32836 31628 32842
rect 31576 32778 31628 32784
rect 31760 32768 31812 32774
rect 31760 32710 31812 32716
rect 31116 32496 31168 32502
rect 31668 32496 31720 32502
rect 31116 32438 31168 32444
rect 31666 32464 31668 32473
rect 31720 32464 31722 32473
rect 31128 31822 31156 32438
rect 31666 32399 31722 32408
rect 31772 32366 31800 32710
rect 31864 32502 31892 33050
rect 31944 32972 31996 32978
rect 31944 32914 31996 32920
rect 31956 32881 31984 32914
rect 32048 32910 32076 33254
rect 32036 32904 32088 32910
rect 31942 32872 31998 32881
rect 32036 32846 32088 32852
rect 31942 32807 31998 32816
rect 31852 32496 31904 32502
rect 31852 32438 31904 32444
rect 31760 32360 31812 32366
rect 31760 32302 31812 32308
rect 31482 32056 31538 32065
rect 31482 31991 31538 32000
rect 31576 32020 31628 32026
rect 31116 31816 31168 31822
rect 31116 31758 31168 31764
rect 31036 31368 31156 31396
rect 30932 31272 30984 31278
rect 30932 31214 30984 31220
rect 30944 30734 30972 31214
rect 31128 31210 31156 31368
rect 31496 31346 31524 31991
rect 31576 31962 31628 31968
rect 31588 31754 31616 31962
rect 31668 31816 31720 31822
rect 31668 31758 31720 31764
rect 31576 31748 31628 31754
rect 31576 31690 31628 31696
rect 31484 31340 31536 31346
rect 31484 31282 31536 31288
rect 31496 31226 31524 31282
rect 31116 31204 31168 31210
rect 31116 31146 31168 31152
rect 31220 31198 31524 31226
rect 30932 30728 30984 30734
rect 30932 30670 30984 30676
rect 30840 30320 30892 30326
rect 30840 30262 30892 30268
rect 31024 29776 31076 29782
rect 31024 29718 31076 29724
rect 30656 29572 30708 29578
rect 30656 29514 30708 29520
rect 30668 29084 30696 29514
rect 31036 29306 31064 29718
rect 31024 29300 31076 29306
rect 31024 29242 31076 29248
rect 30378 29064 30434 29073
rect 30378 28999 30434 29008
rect 30484 29056 30696 29084
rect 30196 28416 30248 28422
rect 30196 28358 30248 28364
rect 30392 28082 30420 28999
rect 30484 28762 30512 29056
rect 30564 28960 30616 28966
rect 30932 28960 30984 28966
rect 30564 28902 30616 28908
rect 30852 28908 30932 28914
rect 30852 28902 30984 28908
rect 30472 28756 30524 28762
rect 30472 28698 30524 28704
rect 30576 28626 30604 28902
rect 30852 28886 30972 28902
rect 30852 28694 30880 28886
rect 31036 28762 31064 29242
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 30840 28688 30892 28694
rect 30840 28630 30892 28636
rect 30564 28620 30616 28626
rect 30564 28562 30616 28568
rect 30656 28552 30708 28558
rect 30656 28494 30708 28500
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 31024 28552 31076 28558
rect 31024 28494 31076 28500
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 29092 28008 29144 28014
rect 29092 27950 29144 27956
rect 30012 28008 30064 28014
rect 30012 27950 30064 27956
rect 28828 27390 28948 27418
rect 28724 26444 28776 26450
rect 28724 26386 28776 26392
rect 28828 25906 28856 27390
rect 29104 27334 29132 27950
rect 29736 27396 29788 27402
rect 29736 27338 29788 27344
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 28908 27124 28960 27130
rect 28908 27066 28960 27072
rect 28920 26314 28948 27066
rect 29564 27062 29592 27270
rect 29552 27056 29604 27062
rect 29552 26998 29604 27004
rect 29748 26994 29776 27338
rect 29644 26988 29696 26994
rect 29644 26930 29696 26936
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 28908 26308 28960 26314
rect 28908 26250 28960 26256
rect 28816 25900 28868 25906
rect 28816 25842 28868 25848
rect 28828 25498 28856 25842
rect 28920 25838 28948 26250
rect 28908 25832 28960 25838
rect 28908 25774 28960 25780
rect 29656 25498 29684 26930
rect 28816 25492 28868 25498
rect 28816 25434 28868 25440
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 28724 25152 28776 25158
rect 28724 25094 28776 25100
rect 28736 24954 28764 25094
rect 28724 24948 28776 24954
rect 28724 24890 28776 24896
rect 29748 24818 29776 26930
rect 30024 26926 30052 27950
rect 30668 27946 30696 28494
rect 30760 28218 30788 28494
rect 30748 28212 30800 28218
rect 30748 28154 30800 28160
rect 30656 27940 30708 27946
rect 30656 27882 30708 27888
rect 30380 27396 30432 27402
rect 30380 27338 30432 27344
rect 30392 27062 30420 27338
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 30380 27056 30432 27062
rect 30380 26998 30432 27004
rect 30196 26988 30248 26994
rect 30196 26930 30248 26936
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 29828 26784 29880 26790
rect 29828 26726 29880 26732
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 28644 24126 28764 24154
rect 28446 23216 28502 23225
rect 28446 23151 28502 23160
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 26516 22976 26568 22982
rect 26516 22918 26568 22924
rect 26148 22034 26200 22040
rect 26252 22066 26372 22094
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25412 21412 25464 21418
rect 25412 21354 25464 21360
rect 25516 21010 25544 21966
rect 25780 21480 25832 21486
rect 25780 21422 25832 21428
rect 25872 21480 25924 21486
rect 25872 21422 25924 21428
rect 25504 21004 25556 21010
rect 25504 20946 25556 20952
rect 25792 20874 25820 21422
rect 25780 20868 25832 20874
rect 25780 20810 25832 20816
rect 25134 20360 25190 20369
rect 25134 20295 25136 20304
rect 25188 20295 25190 20304
rect 25136 20266 25188 20272
rect 25148 19854 25176 20266
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24768 19236 24820 19242
rect 24768 19178 24820 19184
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24596 16590 24624 16934
rect 24780 16590 24808 19178
rect 24872 17814 24900 19314
rect 24964 18426 24992 19790
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24860 17808 24912 17814
rect 24860 17750 24912 17756
rect 24964 17678 24992 18022
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 25056 17202 25084 19450
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25424 19174 25452 19314
rect 25700 19242 25728 20198
rect 25688 19236 25740 19242
rect 25688 19178 25740 19184
rect 25412 19168 25464 19174
rect 25412 19110 25464 19116
rect 25424 18766 25452 19110
rect 25412 18760 25464 18766
rect 25792 18748 25820 20810
rect 25884 19242 25912 21422
rect 26160 21350 26188 22034
rect 26252 21894 26280 22066
rect 26528 21962 26556 22918
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 26160 20942 26188 21286
rect 26344 21146 26372 21898
rect 26884 21616 26936 21622
rect 26528 21554 26740 21570
rect 26884 21558 26936 21564
rect 26976 21616 27028 21622
rect 26976 21558 27028 21564
rect 26528 21548 26752 21554
rect 26528 21542 26700 21548
rect 26528 21486 26556 21542
rect 26700 21490 26752 21496
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 26252 21026 26280 21082
rect 26436 21026 26464 21354
rect 26252 20998 26464 21026
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26146 20360 26202 20369
rect 26146 20295 26202 20304
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 25884 18902 25912 19178
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 25872 18896 25924 18902
rect 25872 18838 25924 18844
rect 25792 18720 25912 18748
rect 25412 18702 25464 18708
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25240 18154 25268 18566
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 25228 18148 25280 18154
rect 25228 18090 25280 18096
rect 25148 17814 25176 18090
rect 25136 17808 25188 17814
rect 25136 17750 25188 17756
rect 25884 17202 25912 18720
rect 25976 18426 26004 19110
rect 26068 18698 26096 19246
rect 26160 18698 26188 20295
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26056 18692 26108 18698
rect 26056 18634 26108 18640
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 25964 18420 26016 18426
rect 25964 18362 26016 18368
rect 26068 18086 26096 18634
rect 26148 18352 26200 18358
rect 26148 18294 26200 18300
rect 26056 18080 26108 18086
rect 26056 18022 26108 18028
rect 26068 17882 26096 18022
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 24214 16144 24270 16153
rect 24136 16102 24214 16130
rect 24214 16079 24216 16088
rect 24268 16079 24270 16088
rect 24216 16050 24268 16056
rect 24504 16046 24532 16458
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 23492 12306 23520 12582
rect 23662 12336 23718 12345
rect 23480 12300 23532 12306
rect 23662 12271 23718 12280
rect 23480 12242 23532 12248
rect 23572 12164 23624 12170
rect 23572 12106 23624 12112
rect 23584 11150 23612 12106
rect 23572 11144 23624 11150
rect 23676 11121 23704 12271
rect 24136 11694 24164 12582
rect 24228 12442 24256 12786
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 24124 11280 24176 11286
rect 24124 11222 24176 11228
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23572 11086 23624 11092
rect 23662 11112 23718 11121
rect 23662 11047 23718 11056
rect 23676 11014 23704 11047
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23204 10736 23256 10742
rect 23204 10678 23256 10684
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23124 8566 23152 9046
rect 23216 8566 23244 10678
rect 23400 10674 23428 10950
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23400 10538 23428 10610
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23400 9654 23428 9862
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23492 9518 23520 9998
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 22940 7534 23060 7562
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22756 7002 22784 7278
rect 22940 7274 22968 7534
rect 23216 7410 23244 8502
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23308 7410 23336 8434
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23492 7818 23520 8230
rect 23388 7812 23440 7818
rect 23388 7754 23440 7760
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23020 7404 23072 7410
rect 23204 7404 23256 7410
rect 23020 7346 23072 7352
rect 23124 7364 23204 7392
rect 22928 7268 22980 7274
rect 22928 7210 22980 7216
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 23032 6644 23060 7346
rect 23124 6798 23152 7364
rect 23204 7346 23256 7352
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23216 6866 23244 7142
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23112 6792 23164 6798
rect 23164 6740 23244 6746
rect 23112 6734 23244 6740
rect 23124 6718 23244 6734
rect 23308 6730 23336 7346
rect 23400 6798 23428 7754
rect 23584 7546 23612 10202
rect 23676 9382 23704 10610
rect 23768 9450 23796 11154
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23860 9926 23888 11018
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23860 8430 23888 9862
rect 23952 8634 23980 10678
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23662 7304 23718 7313
rect 23662 7239 23718 7248
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23112 6656 23164 6662
rect 23032 6616 23112 6644
rect 23032 5710 23060 6616
rect 23112 6598 23164 6604
rect 23112 6180 23164 6186
rect 23112 6122 23164 6128
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 22100 4548 22152 4554
rect 22100 4490 22152 4496
rect 22112 4282 22140 4490
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22204 4078 22232 4966
rect 22388 4146 22416 4966
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 23032 4078 23060 5646
rect 23124 5574 23152 6122
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23124 5302 23152 5510
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23216 5166 23244 6718
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 23216 4826 23244 5102
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23308 4758 23336 6666
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23112 4548 23164 4554
rect 23112 4490 23164 4496
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 21640 4004 21692 4010
rect 21640 3946 21692 3952
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22388 3602 22416 3878
rect 23124 3738 23152 4490
rect 23400 4162 23428 4558
rect 23216 4146 23428 4162
rect 23204 4140 23428 4146
rect 23256 4134 23428 4140
rect 23204 4082 23256 4088
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 23400 3534 23428 4134
rect 23492 4078 23520 6054
rect 23584 5778 23612 6394
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23584 5302 23612 5714
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23676 5030 23704 7239
rect 23768 6322 23796 8298
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7274 23888 7686
rect 23848 7268 23900 7274
rect 23848 7210 23900 7216
rect 23952 7154 23980 8570
rect 24044 8294 24072 11086
rect 24136 10849 24164 11222
rect 24320 11150 24348 13126
rect 24504 12434 24532 15982
rect 24780 13734 24808 16526
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24872 16182 24900 16390
rect 25056 16182 25084 17138
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 24860 16176 24912 16182
rect 24860 16118 24912 16124
rect 25044 16176 25096 16182
rect 25044 16118 25096 16124
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24964 15502 24992 16050
rect 25056 15570 25084 16118
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 24872 14550 24900 14962
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24964 13326 24992 15438
rect 25056 15162 25084 15506
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25056 14498 25084 15098
rect 25228 14884 25280 14890
rect 25228 14826 25280 14832
rect 25320 14884 25372 14890
rect 25320 14826 25372 14832
rect 25056 14482 25176 14498
rect 25056 14476 25188 14482
rect 25056 14470 25136 14476
rect 25056 14074 25084 14470
rect 25136 14418 25188 14424
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 12918 24808 13126
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 24412 12406 24532 12434
rect 24308 11144 24360 11150
rect 24228 11092 24308 11098
rect 24228 11086 24360 11092
rect 24228 11070 24348 11086
rect 24122 10840 24178 10849
rect 24122 10775 24178 10784
rect 24136 10742 24164 10775
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 24124 10532 24176 10538
rect 24124 10474 24176 10480
rect 24136 9586 24164 10474
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24136 7342 24164 9386
rect 24124 7336 24176 7342
rect 24228 7313 24256 11070
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24320 10742 24348 10950
rect 24308 10736 24360 10742
rect 24308 10678 24360 10684
rect 24412 9058 24440 12406
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24780 12102 24808 12174
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24676 11824 24728 11830
rect 24676 11766 24728 11772
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11218 24624 11494
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24596 10674 24624 11154
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24688 10606 24716 11766
rect 24780 11286 24808 12038
rect 25240 11286 25268 14826
rect 25332 14074 25360 14826
rect 25424 14618 25452 16526
rect 25516 16454 25544 17138
rect 25700 16794 25728 17138
rect 25884 17066 25912 17138
rect 25872 17060 25924 17066
rect 25872 17002 25924 17008
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 26160 16674 26188 18294
rect 26252 17814 26280 18906
rect 26344 18834 26372 20742
rect 26528 20398 26556 21422
rect 26896 21010 26924 21558
rect 26884 21004 26936 21010
rect 26884 20946 26936 20952
rect 26792 20800 26844 20806
rect 26792 20742 26844 20748
rect 26804 20602 26832 20742
rect 26792 20596 26844 20602
rect 26792 20538 26844 20544
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 26528 19854 26556 20334
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 26528 19174 26556 19790
rect 26896 19514 26924 20946
rect 26988 20330 27016 21558
rect 26976 20324 27028 20330
rect 26976 20266 27028 20272
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26988 19378 27016 20266
rect 27080 20058 27108 23054
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 27264 22710 27292 22918
rect 27816 22710 27844 22918
rect 27252 22704 27304 22710
rect 27252 22646 27304 22652
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27620 21888 27672 21894
rect 27540 21836 27620 21842
rect 27540 21830 27672 21836
rect 27540 21814 27660 21830
rect 27540 20874 27568 21814
rect 27724 21078 27752 22034
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 27908 21146 27936 21558
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27528 20868 27580 20874
rect 27528 20810 27580 20816
rect 27434 20496 27490 20505
rect 27434 20431 27436 20440
rect 27488 20431 27490 20440
rect 27436 20402 27488 20408
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 27448 19786 27476 20198
rect 27540 20058 27568 20810
rect 27724 20398 27752 21014
rect 27804 20596 27856 20602
rect 27908 20584 27936 21082
rect 27856 20556 27936 20584
rect 27804 20538 27856 20544
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 27804 20392 27856 20398
rect 27908 20369 27936 20402
rect 27804 20334 27856 20340
rect 27894 20360 27950 20369
rect 27816 20210 27844 20334
rect 27894 20295 27950 20304
rect 27724 20182 27844 20210
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27436 19780 27488 19786
rect 27436 19722 27488 19728
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27632 19281 27660 19722
rect 27724 19718 27752 20182
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27618 19272 27674 19281
rect 27618 19207 27674 19216
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26332 18828 26384 18834
rect 26332 18770 26384 18776
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 26424 18420 26476 18426
rect 26424 18362 26476 18368
rect 26332 18216 26384 18222
rect 26332 18158 26384 18164
rect 26344 17882 26372 18158
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26436 17354 26464 18362
rect 26896 18358 26924 18702
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26988 18442 27016 18634
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 26988 18426 27108 18442
rect 26988 18420 27120 18426
rect 26988 18414 27068 18420
rect 26884 18352 26936 18358
rect 26884 18294 26936 18300
rect 26884 17672 26936 17678
rect 26528 17620 26884 17626
rect 26528 17614 26936 17620
rect 26528 17598 26924 17614
rect 26528 17542 26556 17598
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26436 17326 26556 17354
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 26068 16646 26188 16674
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25780 16448 25832 16454
rect 25780 16390 25832 16396
rect 25792 16114 25820 16390
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25516 15570 25544 15846
rect 25504 15564 25556 15570
rect 25504 15506 25556 15512
rect 25884 15162 25912 16594
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25516 13258 25544 13874
rect 25608 13462 25636 14962
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25884 14346 25912 14758
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25596 13456 25648 13462
rect 25596 13398 25648 13404
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25608 12850 25636 13398
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25320 12776 25372 12782
rect 25320 12718 25372 12724
rect 25504 12776 25556 12782
rect 25504 12718 25556 12724
rect 25332 12220 25360 12718
rect 25412 12232 25464 12238
rect 25332 12192 25412 12220
rect 25412 12174 25464 12180
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 25228 11280 25280 11286
rect 25228 11222 25280 11228
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 24952 11076 25004 11082
rect 24952 11018 25004 11024
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24964 10538 24992 11018
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 25240 10470 25268 10610
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25240 9722 25268 9930
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25332 9586 25360 11154
rect 25424 11014 25452 12174
rect 25516 11642 25544 12718
rect 25608 12442 25636 12786
rect 25700 12714 25728 13126
rect 25792 12850 25820 13262
rect 26068 13190 26096 16646
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26160 13938 26188 16526
rect 26424 15360 26476 15366
rect 26424 15302 26476 15308
rect 26436 15026 26464 15302
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26252 13530 26280 13874
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26528 13462 26556 17326
rect 26712 16998 26740 17478
rect 26700 16992 26752 16998
rect 26700 16934 26752 16940
rect 26712 16114 26740 16934
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26712 15638 26740 16050
rect 26700 15632 26752 15638
rect 26700 15574 26752 15580
rect 26712 14958 26740 15574
rect 26896 15366 26924 17598
rect 26988 16658 27016 18414
rect 27068 18362 27120 18368
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27264 18057 27292 18226
rect 27250 18048 27306 18057
rect 27080 18006 27250 18034
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 27080 16153 27108 18006
rect 27250 17983 27306 17992
rect 27632 17746 27660 18566
rect 27724 18222 27752 19654
rect 28000 19514 28028 21966
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28080 20868 28132 20874
rect 28080 20810 28132 20816
rect 27988 19508 28040 19514
rect 27988 19450 28040 19456
rect 28000 18970 28028 19450
rect 28092 19310 28120 20810
rect 28184 20602 28212 21082
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28264 20528 28316 20534
rect 28262 20496 28264 20505
rect 28316 20496 28318 20505
rect 28262 20431 28318 20440
rect 28368 20398 28396 21966
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28644 21486 28672 21558
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 28552 21146 28580 21422
rect 28540 21140 28592 21146
rect 28540 21082 28592 21088
rect 28736 21026 28764 24126
rect 29564 23186 29592 24210
rect 29840 24138 29868 26726
rect 29920 26444 29972 26450
rect 30024 26432 30052 26862
rect 30104 26444 30156 26450
rect 30024 26404 30104 26432
rect 29920 26386 29972 26392
rect 30104 26386 30156 26392
rect 29932 25906 29960 26386
rect 30208 25906 30236 26930
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 30300 26382 30328 26862
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 29920 25900 29972 25906
rect 29920 25842 29972 25848
rect 30196 25900 30248 25906
rect 30196 25842 30248 25848
rect 29932 25362 29960 25842
rect 30012 25832 30064 25838
rect 30012 25774 30064 25780
rect 29920 25356 29972 25362
rect 29920 25298 29972 25304
rect 30024 25294 30052 25774
rect 30208 25378 30236 25842
rect 30392 25838 30420 26998
rect 30576 26382 30604 27270
rect 30668 26790 30696 27882
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 30748 27600 30800 27606
rect 30748 27542 30800 27548
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30472 26308 30524 26314
rect 30472 26250 30524 26256
rect 30380 25832 30432 25838
rect 30380 25774 30432 25780
rect 30208 25350 30420 25378
rect 30012 25288 30064 25294
rect 30012 25230 30064 25236
rect 30208 24954 30236 25350
rect 30288 25288 30340 25294
rect 30288 25230 30340 25236
rect 30196 24948 30248 24954
rect 30196 24890 30248 24896
rect 30300 24750 30328 25230
rect 30392 24818 30420 25350
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30288 24744 30340 24750
rect 30288 24686 30340 24692
rect 30300 24274 30328 24686
rect 30484 24682 30512 26250
rect 30564 26240 30616 26246
rect 30564 26182 30616 26188
rect 30576 25362 30604 26182
rect 30760 25974 30788 27542
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30852 26518 30880 26794
rect 30840 26512 30892 26518
rect 30840 26454 30892 26460
rect 30840 26240 30892 26246
rect 30840 26182 30892 26188
rect 30748 25968 30800 25974
rect 30748 25910 30800 25916
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30668 24886 30696 25842
rect 30760 24954 30788 25910
rect 30852 25226 30880 26182
rect 30944 26042 30972 27814
rect 30932 26036 30984 26042
rect 30932 25978 30984 25984
rect 30932 25832 30984 25838
rect 30932 25774 30984 25780
rect 30840 25220 30892 25226
rect 30840 25162 30892 25168
rect 30748 24948 30800 24954
rect 30748 24890 30800 24896
rect 30656 24880 30708 24886
rect 30656 24822 30708 24828
rect 30472 24676 30524 24682
rect 30472 24618 30524 24624
rect 30288 24268 30340 24274
rect 30288 24210 30340 24216
rect 29828 24132 29880 24138
rect 29828 24074 29880 24080
rect 30668 24070 30696 24822
rect 30944 24818 30972 25774
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 31036 23730 31064 28494
rect 31128 27674 31156 31146
rect 31220 28762 31248 31198
rect 31484 30320 31536 30326
rect 31484 30262 31536 30268
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31404 29510 31432 29990
rect 31496 29714 31524 30262
rect 31484 29708 31536 29714
rect 31484 29650 31536 29656
rect 31392 29504 31444 29510
rect 31392 29446 31444 29452
rect 31404 29170 31432 29446
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31496 28966 31524 29650
rect 31484 28960 31536 28966
rect 31484 28902 31536 28908
rect 31588 28762 31616 31690
rect 31680 30122 31708 31758
rect 31772 31482 31800 32302
rect 31956 32298 31984 32807
rect 32048 32570 32076 32846
rect 32036 32564 32088 32570
rect 32036 32506 32088 32512
rect 31944 32292 31996 32298
rect 31944 32234 31996 32240
rect 31956 31822 31984 32234
rect 32140 31958 32168 33458
rect 32128 31952 32180 31958
rect 32128 31894 32180 31900
rect 31944 31816 31996 31822
rect 31944 31758 31996 31764
rect 32232 31754 32260 35634
rect 32416 35290 32444 36654
rect 32600 35834 32628 36654
rect 34808 36378 34836 37130
rect 34900 36786 34928 37334
rect 36740 37330 36768 37431
rect 36728 37324 36780 37330
rect 36728 37266 36780 37272
rect 36544 37188 36596 37194
rect 36544 37130 36596 37136
rect 35900 37120 35952 37126
rect 35900 37062 35952 37068
rect 34888 36780 34940 36786
rect 34888 36722 34940 36728
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34796 36372 34848 36378
rect 34796 36314 34848 36320
rect 34612 36168 34664 36174
rect 34612 36110 34664 36116
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 35806 36136 35862 36145
rect 32588 35828 32640 35834
rect 32588 35770 32640 35776
rect 34624 35698 34652 36110
rect 32588 35692 32640 35698
rect 32588 35634 32640 35640
rect 34612 35692 34664 35698
rect 34612 35634 34664 35640
rect 32404 35284 32456 35290
rect 32404 35226 32456 35232
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 32416 34066 32444 34546
rect 32404 34060 32456 34066
rect 32404 34002 32456 34008
rect 32312 33924 32364 33930
rect 32312 33866 32364 33872
rect 32324 32570 32352 33866
rect 32416 33522 32444 34002
rect 32404 33516 32456 33522
rect 32404 33458 32456 33464
rect 32496 32972 32548 32978
rect 32496 32914 32548 32920
rect 32404 32768 32456 32774
rect 32404 32710 32456 32716
rect 32312 32564 32364 32570
rect 32312 32506 32364 32512
rect 32416 32434 32444 32710
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32312 32360 32364 32366
rect 32312 32302 32364 32308
rect 32140 31726 32260 31754
rect 31760 31476 31812 31482
rect 31760 31418 31812 31424
rect 32036 30592 32088 30598
rect 32036 30534 32088 30540
rect 31852 30388 31904 30394
rect 31852 30330 31904 30336
rect 31668 30116 31720 30122
rect 31668 30058 31720 30064
rect 31680 29646 31708 30058
rect 31760 30048 31812 30054
rect 31760 29990 31812 29996
rect 31668 29640 31720 29646
rect 31668 29582 31720 29588
rect 31772 29170 31800 29990
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31576 28756 31628 28762
rect 31576 28698 31628 28704
rect 31668 28756 31720 28762
rect 31668 28698 31720 28704
rect 31576 28620 31628 28626
rect 31576 28562 31628 28568
rect 31392 28076 31444 28082
rect 31392 28018 31444 28024
rect 31484 28076 31536 28082
rect 31484 28018 31536 28024
rect 31116 27668 31168 27674
rect 31116 27610 31168 27616
rect 31116 27532 31168 27538
rect 31116 27474 31168 27480
rect 31128 26994 31156 27474
rect 31208 27464 31260 27470
rect 31208 27406 31260 27412
rect 31116 26988 31168 26994
rect 31116 26930 31168 26936
rect 31220 26858 31248 27406
rect 31300 27124 31352 27130
rect 31300 27066 31352 27072
rect 31208 26852 31260 26858
rect 31208 26794 31260 26800
rect 31208 26036 31260 26042
rect 31208 25978 31260 25984
rect 31220 25158 31248 25978
rect 31312 25906 31340 27066
rect 31404 25974 31432 28018
rect 31496 27878 31524 28018
rect 31588 27946 31616 28562
rect 31680 28014 31708 28698
rect 31668 28008 31720 28014
rect 31668 27950 31720 27956
rect 31576 27940 31628 27946
rect 31576 27882 31628 27888
rect 31484 27872 31536 27878
rect 31484 27814 31536 27820
rect 31496 27674 31524 27814
rect 31484 27668 31536 27674
rect 31484 27610 31536 27616
rect 31484 26988 31536 26994
rect 31484 26930 31536 26936
rect 31496 26790 31524 26930
rect 31576 26920 31628 26926
rect 31576 26862 31628 26868
rect 31484 26784 31536 26790
rect 31484 26726 31536 26732
rect 31496 26382 31524 26726
rect 31484 26376 31536 26382
rect 31484 26318 31536 26324
rect 31392 25968 31444 25974
rect 31392 25910 31444 25916
rect 31588 25906 31616 26862
rect 31300 25900 31352 25906
rect 31300 25842 31352 25848
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 31208 25152 31260 25158
rect 31208 25094 31260 25100
rect 31116 24948 31168 24954
rect 31116 24890 31168 24896
rect 31128 24818 31156 24890
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 30840 23248 30892 23254
rect 30840 23190 30892 23196
rect 29552 23180 29604 23186
rect 29552 23122 29604 23128
rect 29460 23044 29512 23050
rect 29460 22986 29512 22992
rect 29472 22778 29500 22986
rect 29460 22772 29512 22778
rect 29460 22714 29512 22720
rect 29276 22636 29328 22642
rect 29276 22578 29328 22584
rect 29000 22432 29052 22438
rect 29000 22374 29052 22380
rect 28908 21888 28960 21894
rect 28908 21830 28960 21836
rect 28552 20998 28764 21026
rect 28920 21010 28948 21830
rect 28908 21004 28960 21010
rect 28356 20392 28408 20398
rect 28262 20360 28318 20369
rect 28356 20334 28408 20340
rect 28262 20295 28318 20304
rect 28276 19378 28304 20295
rect 28368 19922 28396 20334
rect 28356 19916 28408 19922
rect 28356 19858 28408 19864
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28460 19514 28488 19790
rect 28448 19508 28500 19514
rect 28448 19450 28500 19456
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28552 19334 28580 20998
rect 28908 20946 28960 20952
rect 28908 20868 28960 20874
rect 28908 20810 28960 20816
rect 28920 20466 28948 20810
rect 29012 20534 29040 22374
rect 29092 22024 29144 22030
rect 29092 21966 29144 21972
rect 29104 20874 29132 21966
rect 29092 20868 29144 20874
rect 29092 20810 29144 20816
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 29000 20392 29052 20398
rect 28906 20360 28962 20369
rect 28962 20340 29000 20346
rect 28962 20334 29052 20340
rect 28962 20318 29040 20334
rect 28906 20295 28962 20304
rect 28816 20256 28868 20262
rect 28868 20216 28948 20244
rect 28816 20198 28868 20204
rect 28920 20058 28948 20216
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 28906 19952 28962 19961
rect 28906 19887 28908 19896
rect 28960 19887 28962 19896
rect 28908 19858 28960 19864
rect 29104 19666 29132 20810
rect 29184 20324 29236 20330
rect 29184 20266 29236 20272
rect 28920 19638 29132 19666
rect 28920 19514 28948 19638
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 29196 19378 29224 20266
rect 29184 19372 29236 19378
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 28460 19242 28488 19314
rect 28552 19306 28764 19334
rect 29184 19314 29236 19320
rect 28448 19236 28500 19242
rect 28448 19178 28500 19184
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 28264 18692 28316 18698
rect 28264 18634 28316 18640
rect 28276 18290 28304 18634
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27160 17536 27212 17542
rect 27160 17478 27212 17484
rect 27172 17338 27200 17478
rect 27540 17338 27568 17614
rect 27724 17610 27752 18158
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27620 17332 27672 17338
rect 27620 17274 27672 17280
rect 27252 17264 27304 17270
rect 27252 17206 27304 17212
rect 27436 17264 27488 17270
rect 27632 17218 27660 17274
rect 27436 17206 27488 17212
rect 27264 16697 27292 17206
rect 27250 16688 27306 16697
rect 27250 16623 27306 16632
rect 27066 16144 27122 16153
rect 27264 16114 27292 16623
rect 27066 16079 27122 16088
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27252 16108 27304 16114
rect 27252 16050 27304 16056
rect 26884 15360 26936 15366
rect 26884 15302 26936 15308
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26700 14000 26752 14006
rect 26700 13942 26752 13948
rect 26516 13456 26568 13462
rect 26516 13398 26568 13404
rect 26056 13184 26108 13190
rect 26056 13126 26108 13132
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25688 12708 25740 12714
rect 25688 12650 25740 12656
rect 25792 12646 25820 12786
rect 25780 12640 25832 12646
rect 25780 12582 25832 12588
rect 25964 12640 26016 12646
rect 25964 12582 26016 12588
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25792 11898 25820 12582
rect 25976 12306 26004 12582
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 26344 12238 26372 13126
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 26344 11830 26372 12174
rect 26332 11824 26384 11830
rect 26332 11766 26384 11772
rect 25596 11688 25648 11694
rect 25516 11636 25596 11642
rect 25516 11630 25648 11636
rect 25516 11614 25636 11630
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25424 10742 25452 10950
rect 25412 10736 25464 10742
rect 25412 10678 25464 10684
rect 25608 10674 25636 11614
rect 26240 11620 26292 11626
rect 26240 11562 26292 11568
rect 26056 11212 26108 11218
rect 26056 11154 26108 11160
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25976 10810 26004 11086
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24688 9110 24716 9454
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 9178 25084 9318
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 24320 9030 24440 9058
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24492 9036 24544 9042
rect 24320 8362 24348 9030
rect 24492 8978 24544 8984
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 24308 8356 24360 8362
rect 24308 8298 24360 8304
rect 24412 7886 24440 8774
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24504 7410 24532 8978
rect 24766 8936 24822 8945
rect 24766 8871 24768 8880
rect 24820 8871 24822 8880
rect 24768 8842 24820 8848
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24688 8634 24716 8774
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24780 8294 24808 8434
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24124 7278 24176 7284
rect 24214 7304 24270 7313
rect 24214 7239 24270 7248
rect 24780 7206 24808 7686
rect 24872 7410 24900 8570
rect 25056 8566 25084 8978
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25148 8634 25176 8910
rect 25608 8809 25636 8978
rect 25594 8800 25650 8809
rect 25594 8735 25650 8744
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 25148 8498 25176 8570
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25056 7818 25084 8026
rect 25148 7886 25176 8434
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25044 7812 25096 7818
rect 25044 7754 25096 7760
rect 25056 7546 25084 7754
rect 25240 7750 25268 8366
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25332 7818 25360 8230
rect 25504 8016 25556 8022
rect 25504 7958 25556 7964
rect 25320 7812 25372 7818
rect 25320 7754 25372 7760
rect 25228 7744 25280 7750
rect 25228 7686 25280 7692
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 24768 7200 24820 7206
rect 23952 7126 24072 7154
rect 24768 7142 24820 7148
rect 24044 6458 24072 7126
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 23860 5710 23888 6054
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23952 5370 23980 6326
rect 24688 6254 24716 6734
rect 24780 6322 24808 7142
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 25056 6458 25084 6734
rect 25148 6458 25176 7346
rect 25240 6798 25268 7686
rect 25332 7274 25360 7754
rect 25320 7268 25372 7274
rect 25320 7210 25372 7216
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24688 5370 24716 6190
rect 25240 5710 25268 6598
rect 25332 6322 25360 7210
rect 25516 6866 25544 7958
rect 25700 7886 25728 9590
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25780 9104 25832 9110
rect 25780 9046 25832 9052
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25792 7410 25820 9046
rect 25884 8362 25912 9522
rect 25976 9518 26004 9590
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 26068 9466 26096 11154
rect 26148 10532 26200 10538
rect 26148 10474 26200 10480
rect 26160 9674 26188 10474
rect 26252 10470 26280 11562
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 26252 10130 26280 10406
rect 26332 10192 26384 10198
rect 26332 10134 26384 10140
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26160 9646 26280 9674
rect 26252 9518 26280 9646
rect 26148 9512 26200 9518
rect 26068 9460 26148 9466
rect 26068 9454 26200 9460
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 25872 8356 25924 8362
rect 25872 8298 25924 8304
rect 25884 8022 25912 8298
rect 25872 8016 25924 8022
rect 25872 7958 25924 7964
rect 25976 7868 26004 9454
rect 26068 9438 26188 9454
rect 26068 9110 26096 9438
rect 26056 9104 26108 9110
rect 26056 9046 26108 9052
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 26146 8936 26202 8945
rect 26068 8090 26096 8910
rect 26252 8922 26280 9454
rect 26202 8894 26280 8922
rect 26146 8871 26202 8880
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26056 7880 26108 7886
rect 25976 7840 26056 7868
rect 26056 7822 26108 7828
rect 26160 7410 26188 8871
rect 26240 8832 26292 8838
rect 26344 8820 26372 10134
rect 26436 9586 26464 12922
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26620 11626 26648 12174
rect 26608 11620 26660 11626
rect 26608 11562 26660 11568
rect 26712 11354 26740 13942
rect 26884 13456 26936 13462
rect 26884 13398 26936 13404
rect 26896 13326 26924 13398
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26988 12918 27016 15030
rect 27172 13734 27200 16050
rect 27448 15978 27476 17206
rect 27540 17190 27660 17218
rect 27540 16726 27568 17190
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27528 16720 27580 16726
rect 27528 16662 27580 16668
rect 27528 16584 27580 16590
rect 27632 16538 27660 17070
rect 27724 16726 27752 17546
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27712 16720 27764 16726
rect 27712 16662 27764 16668
rect 27580 16532 27660 16538
rect 27528 16526 27660 16532
rect 27540 16510 27660 16526
rect 27632 16250 27660 16510
rect 27712 16516 27764 16522
rect 27712 16458 27764 16464
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27620 16108 27672 16114
rect 27724 16096 27752 16458
rect 27672 16068 27752 16096
rect 27620 16050 27672 16056
rect 27436 15972 27488 15978
rect 27436 15914 27488 15920
rect 27816 15502 27844 16730
rect 28092 16726 28120 18022
rect 28276 17610 28304 18226
rect 28460 18086 28488 19178
rect 28540 18896 28592 18902
rect 28540 18838 28592 18844
rect 28448 18080 28500 18086
rect 28448 18022 28500 18028
rect 28264 17604 28316 17610
rect 28264 17546 28316 17552
rect 28276 17202 28304 17546
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 27896 16720 27948 16726
rect 27896 16662 27948 16668
rect 28080 16720 28132 16726
rect 28080 16662 28132 16668
rect 27804 15496 27856 15502
rect 27804 15438 27856 15444
rect 27908 15450 27936 16662
rect 28092 16454 28120 16662
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28080 16176 28132 16182
rect 28080 16118 28132 16124
rect 27988 15904 28040 15910
rect 27988 15846 28040 15852
rect 28000 15570 28028 15846
rect 28092 15706 28120 16118
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 27988 15564 28040 15570
rect 27988 15506 28040 15512
rect 28276 15502 28304 16390
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28368 15706 28396 15846
rect 28356 15700 28408 15706
rect 28356 15642 28408 15648
rect 28264 15496 28316 15502
rect 27816 14958 27844 15438
rect 27908 15422 28028 15450
rect 28264 15438 28316 15444
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27804 14952 27856 14958
rect 27804 14894 27856 14900
rect 27436 14340 27488 14346
rect 27436 14282 27488 14288
rect 27344 14000 27396 14006
rect 27344 13942 27396 13948
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 26976 12912 27028 12918
rect 26976 12854 27028 12860
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26804 11898 26832 12786
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26514 10024 26570 10033
rect 26514 9959 26570 9968
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 26436 9042 26464 9522
rect 26528 9518 26556 9959
rect 26712 9926 26740 11086
rect 26988 10742 27016 12854
rect 27080 11150 27108 13126
rect 27356 12345 27384 13942
rect 27342 12336 27398 12345
rect 27342 12271 27398 12280
rect 27448 11354 27476 14282
rect 27816 13326 27844 14894
rect 27908 14074 27936 14962
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 28000 13734 28028 15422
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 28552 13530 28580 18838
rect 28736 17746 28764 19306
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 29104 18766 29132 19246
rect 29288 18970 29316 22578
rect 29564 22166 29592 23122
rect 30380 23044 30432 23050
rect 30380 22986 30432 22992
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 30116 22438 30144 22578
rect 30012 22432 30064 22438
rect 30012 22374 30064 22380
rect 30104 22432 30156 22438
rect 30104 22374 30156 22380
rect 29552 22160 29604 22166
rect 29552 22102 29604 22108
rect 30024 21622 30052 22374
rect 30116 22030 30144 22374
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30392 21962 30420 22986
rect 30852 22642 30880 23190
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30380 21956 30432 21962
rect 30380 21898 30432 21904
rect 30484 21690 30512 22578
rect 31116 22092 31168 22098
rect 31116 22034 31168 22040
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30472 21684 30524 21690
rect 30472 21626 30524 21632
rect 30012 21616 30064 21622
rect 30012 21558 30064 21564
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 29920 21480 29972 21486
rect 29920 21422 29972 21428
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29748 20942 29776 21286
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29736 20324 29788 20330
rect 29736 20266 29788 20272
rect 29644 19916 29696 19922
rect 29644 19858 29696 19864
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29276 18964 29328 18970
rect 29276 18906 29328 18912
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 29564 18698 29592 19790
rect 29656 19514 29684 19858
rect 29748 19854 29776 20266
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29828 19780 29880 19786
rect 29828 19722 29880 19728
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 29840 19378 29868 19722
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29552 18692 29604 18698
rect 29552 18634 29604 18640
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 28724 17740 28776 17746
rect 28724 17682 28776 17688
rect 28630 16688 28686 16697
rect 28630 16623 28632 16632
rect 28684 16623 28686 16632
rect 28632 16594 28684 16600
rect 29012 15094 29040 18566
rect 29932 17882 29960 21422
rect 30012 21140 30064 21146
rect 30012 21082 30064 21088
rect 30024 20534 30052 21082
rect 30012 20528 30064 20534
rect 30012 20470 30064 20476
rect 30668 20262 30696 21490
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 30116 19378 30144 19994
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 30392 19242 30420 19450
rect 30576 19310 30604 19790
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30564 19304 30616 19310
rect 30564 19246 30616 19252
rect 30380 19236 30432 19242
rect 30380 19178 30432 19184
rect 30196 19168 30248 19174
rect 30196 19110 30248 19116
rect 30104 18896 30156 18902
rect 30010 18864 30066 18873
rect 30104 18838 30156 18844
rect 30010 18799 30066 18808
rect 30024 18766 30052 18799
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 30024 18630 30052 18702
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 30116 18578 30144 18838
rect 30208 18766 30236 19110
rect 30288 18896 30340 18902
rect 30288 18838 30340 18844
rect 30196 18760 30248 18766
rect 30196 18702 30248 18708
rect 30300 18578 30328 18838
rect 30116 18550 30328 18578
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 30116 17678 30144 18158
rect 29828 17672 29880 17678
rect 29828 17614 29880 17620
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 29644 17060 29696 17066
rect 29644 17002 29696 17008
rect 29656 16794 29684 17002
rect 29644 16788 29696 16794
rect 29644 16730 29696 16736
rect 29368 16720 29420 16726
rect 29368 16662 29420 16668
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29196 15978 29224 16526
rect 29184 15972 29236 15978
rect 29184 15914 29236 15920
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 29092 15020 29144 15026
rect 29196 15008 29224 15914
rect 29380 15162 29408 16662
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 29656 16522 29684 16594
rect 29644 16516 29696 16522
rect 29644 16458 29696 16464
rect 29656 16250 29684 16458
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 29644 16244 29696 16250
rect 29644 16186 29696 16192
rect 29748 15502 29776 16390
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29840 15162 29868 17614
rect 30116 16454 30144 17614
rect 30300 16794 30328 18550
rect 30668 18358 30696 19654
rect 30760 18970 30788 21898
rect 30840 21684 30892 21690
rect 30840 21626 30892 21632
rect 30852 20942 30880 21626
rect 31128 21418 31156 22034
rect 31116 21412 31168 21418
rect 31116 21354 31168 21360
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 30840 20936 30892 20942
rect 30840 20878 30892 20884
rect 30852 20466 30880 20878
rect 30840 20460 30892 20466
rect 30840 20402 30892 20408
rect 30932 20392 30984 20398
rect 30932 20334 30984 20340
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30852 19854 30880 20198
rect 30840 19848 30892 19854
rect 30840 19790 30892 19796
rect 30852 18970 30880 19790
rect 30944 19718 30972 20334
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30748 18964 30800 18970
rect 30748 18906 30800 18912
rect 30840 18964 30892 18970
rect 30840 18906 30892 18912
rect 30944 18680 30972 19654
rect 31036 19514 31064 21286
rect 31128 21078 31156 21354
rect 31116 21072 31168 21078
rect 31116 21014 31168 21020
rect 31128 19922 31156 21014
rect 31116 19916 31168 19922
rect 31116 19858 31168 19864
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 31128 18766 31156 19858
rect 31220 18902 31248 25094
rect 31588 24886 31616 25842
rect 31576 24880 31628 24886
rect 31576 24822 31628 24828
rect 31864 24698 31892 30330
rect 32048 29850 32076 30534
rect 32036 29844 32088 29850
rect 32036 29786 32088 29792
rect 32140 29594 32168 31726
rect 32324 31210 32352 32302
rect 32508 31822 32536 32914
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 32508 31414 32536 31758
rect 32496 31408 32548 31414
rect 32496 31350 32548 31356
rect 32312 31204 32364 31210
rect 32312 31146 32364 31152
rect 32220 30660 32272 30666
rect 32220 30602 32272 30608
rect 32232 30546 32260 30602
rect 32232 30518 32444 30546
rect 32416 30122 32444 30518
rect 32600 30394 32628 35634
rect 33782 34640 33838 34649
rect 33416 34604 33468 34610
rect 34716 34610 34744 36110
rect 35806 36071 35862 36080
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 33782 34575 33838 34584
rect 34704 34604 34756 34610
rect 33416 34546 33468 34552
rect 33324 33924 33376 33930
rect 33324 33866 33376 33872
rect 33336 33658 33364 33866
rect 33324 33652 33376 33658
rect 33324 33594 33376 33600
rect 32956 33312 33008 33318
rect 32956 33254 33008 33260
rect 32772 32904 32824 32910
rect 32770 32872 32772 32881
rect 32824 32872 32826 32881
rect 32968 32842 32996 33254
rect 33428 33017 33456 34546
rect 33796 34542 33824 34575
rect 34704 34546 34756 34552
rect 35820 34542 35848 36071
rect 35912 35766 35940 37062
rect 35900 35760 35952 35766
rect 35900 35702 35952 35708
rect 36556 34678 36584 37130
rect 36832 35494 36860 37590
rect 37200 36786 37228 38791
rect 37280 37256 37332 37262
rect 37280 37198 37332 37204
rect 37188 36780 37240 36786
rect 37188 36722 37240 36728
rect 36728 35488 36780 35494
rect 36728 35430 36780 35436
rect 36820 35488 36872 35494
rect 36820 35430 36872 35436
rect 36740 35290 36768 35430
rect 36728 35284 36780 35290
rect 36728 35226 36780 35232
rect 37188 35148 37240 35154
rect 37188 35090 37240 35096
rect 36728 35080 36780 35086
rect 36728 35022 36780 35028
rect 36544 34672 36596 34678
rect 36544 34614 36596 34620
rect 36740 34610 36768 35022
rect 37200 34785 37228 35090
rect 37186 34776 37242 34785
rect 37186 34711 37242 34720
rect 36728 34604 36780 34610
rect 36728 34546 36780 34552
rect 33784 34536 33836 34542
rect 35808 34536 35860 34542
rect 33836 34496 34008 34524
rect 33784 34478 33836 34484
rect 33600 33108 33652 33114
rect 33600 33050 33652 33056
rect 33414 33008 33470 33017
rect 33414 32943 33470 32952
rect 32770 32807 32826 32816
rect 32956 32836 33008 32842
rect 32956 32778 33008 32784
rect 32864 32496 32916 32502
rect 32864 32438 32916 32444
rect 32876 31482 32904 32438
rect 32968 32434 32996 32778
rect 32956 32428 33008 32434
rect 32956 32370 33008 32376
rect 32968 31890 32996 32370
rect 33232 32360 33284 32366
rect 33232 32302 33284 32308
rect 33416 32360 33468 32366
rect 33416 32302 33468 32308
rect 33244 31890 33272 32302
rect 32956 31884 33008 31890
rect 32956 31826 33008 31832
rect 33232 31884 33284 31890
rect 33232 31826 33284 31832
rect 33244 31754 33272 31826
rect 33244 31726 33364 31754
rect 32864 31476 32916 31482
rect 32864 31418 32916 31424
rect 33048 31136 33100 31142
rect 33048 31078 33100 31084
rect 33060 30666 33088 31078
rect 33048 30660 33100 30666
rect 33048 30602 33100 30608
rect 32588 30388 32640 30394
rect 32588 30330 32640 30336
rect 32404 30116 32456 30122
rect 32404 30058 32456 30064
rect 32588 30116 32640 30122
rect 32588 30058 32640 30064
rect 32048 29566 32168 29594
rect 32048 26042 32076 29566
rect 32128 29504 32180 29510
rect 32128 29446 32180 29452
rect 32312 29504 32364 29510
rect 32312 29446 32364 29452
rect 32140 29322 32168 29446
rect 32140 29306 32260 29322
rect 32140 29300 32272 29306
rect 32140 29294 32220 29300
rect 32140 29170 32168 29294
rect 32220 29242 32272 29248
rect 32324 29170 32352 29446
rect 32128 29164 32180 29170
rect 32128 29106 32180 29112
rect 32312 29164 32364 29170
rect 32312 29106 32364 29112
rect 32140 28218 32168 29106
rect 32324 28558 32352 29106
rect 32312 28552 32364 28558
rect 32312 28494 32364 28500
rect 32128 28212 32180 28218
rect 32128 28154 32180 28160
rect 32128 27328 32180 27334
rect 32128 27270 32180 27276
rect 32140 26382 32168 27270
rect 32416 27062 32444 30058
rect 32600 29510 32628 30058
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32588 29504 32640 29510
rect 32588 29446 32640 29452
rect 32968 29170 32996 29786
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 33244 29238 33272 29582
rect 33232 29232 33284 29238
rect 33232 29174 33284 29180
rect 32956 29164 33008 29170
rect 32956 29106 33008 29112
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 33140 29096 33192 29102
rect 33140 29038 33192 29044
rect 32680 28484 32732 28490
rect 32680 28426 32732 28432
rect 32496 28416 32548 28422
rect 32496 28358 32548 28364
rect 32508 27946 32536 28358
rect 32496 27940 32548 27946
rect 32496 27882 32548 27888
rect 32692 27538 32720 28426
rect 32772 28416 32824 28422
rect 32772 28358 32824 28364
rect 32784 28218 32812 28358
rect 32772 28212 32824 28218
rect 32772 28154 32824 28160
rect 32680 27532 32732 27538
rect 32680 27474 32732 27480
rect 32588 27464 32640 27470
rect 32588 27406 32640 27412
rect 32404 27056 32456 27062
rect 32404 26998 32456 27004
rect 32496 26852 32548 26858
rect 32496 26794 32548 26800
rect 32404 26580 32456 26586
rect 32404 26522 32456 26528
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 32220 26308 32272 26314
rect 32220 26250 32272 26256
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 32036 25832 32088 25838
rect 32036 25774 32088 25780
rect 32048 25498 32076 25774
rect 32232 25498 32260 26250
rect 32036 25492 32088 25498
rect 32036 25434 32088 25440
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32416 24750 32444 26522
rect 32508 26314 32536 26794
rect 32496 26308 32548 26314
rect 32496 26250 32548 26256
rect 32600 25294 32628 27406
rect 32692 27130 32720 27474
rect 32876 27130 32904 29038
rect 33152 28694 33180 29038
rect 33140 28688 33192 28694
rect 33140 28630 33192 28636
rect 32956 28144 33008 28150
rect 32956 28086 33008 28092
rect 32968 27674 32996 28086
rect 33152 28082 33180 28630
rect 33336 28626 33364 31726
rect 33428 30802 33456 32302
rect 33612 31226 33640 33050
rect 33692 32836 33744 32842
rect 33692 32778 33744 32784
rect 33704 31958 33732 32778
rect 33692 31952 33744 31958
rect 33692 31894 33744 31900
rect 33704 31346 33732 31894
rect 33784 31748 33836 31754
rect 33784 31690 33836 31696
rect 33876 31748 33928 31754
rect 33876 31690 33928 31696
rect 33692 31340 33744 31346
rect 33692 31282 33744 31288
rect 33796 31226 33824 31690
rect 33888 31482 33916 31690
rect 33876 31476 33928 31482
rect 33876 31418 33928 31424
rect 33612 31198 33824 31226
rect 33416 30796 33468 30802
rect 33416 30738 33468 30744
rect 33508 30660 33560 30666
rect 33508 30602 33560 30608
rect 33520 29850 33548 30602
rect 33508 29844 33560 29850
rect 33508 29786 33560 29792
rect 33416 29640 33468 29646
rect 33416 29582 33468 29588
rect 33428 28762 33456 29582
rect 33416 28756 33468 28762
rect 33416 28698 33468 28704
rect 33324 28620 33376 28626
rect 33324 28562 33376 28568
rect 33140 28076 33192 28082
rect 33140 28018 33192 28024
rect 33336 28014 33364 28562
rect 33612 28370 33640 31198
rect 33784 30116 33836 30122
rect 33784 30058 33836 30064
rect 33692 29096 33744 29102
rect 33692 29038 33744 29044
rect 33704 28490 33732 29038
rect 33796 28966 33824 30058
rect 33784 28960 33836 28966
rect 33784 28902 33836 28908
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33692 28484 33744 28490
rect 33692 28426 33744 28432
rect 33796 28370 33824 28494
rect 33612 28342 33824 28370
rect 33692 28144 33744 28150
rect 33692 28086 33744 28092
rect 33600 28076 33652 28082
rect 33600 28018 33652 28024
rect 33324 28008 33376 28014
rect 33324 27950 33376 27956
rect 32956 27668 33008 27674
rect 32956 27610 33008 27616
rect 32968 27470 32996 27610
rect 32956 27464 33008 27470
rect 32956 27406 33008 27412
rect 32680 27124 32732 27130
rect 32680 27066 32732 27072
rect 32864 27124 32916 27130
rect 32864 27066 32916 27072
rect 32680 26988 32732 26994
rect 32680 26930 32732 26936
rect 32692 25906 32720 26930
rect 33232 26920 33284 26926
rect 33232 26862 33284 26868
rect 33244 26314 33272 26862
rect 33336 26790 33364 27950
rect 33508 27872 33560 27878
rect 33508 27814 33560 27820
rect 33520 27538 33548 27814
rect 33508 27532 33560 27538
rect 33508 27474 33560 27480
rect 33520 27334 33548 27474
rect 33612 27402 33640 28018
rect 33600 27396 33652 27402
rect 33600 27338 33652 27344
rect 33508 27328 33560 27334
rect 33508 27270 33560 27276
rect 33416 26988 33468 26994
rect 33416 26930 33468 26936
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 33336 26450 33364 26726
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33232 26308 33284 26314
rect 33232 26250 33284 26256
rect 32680 25900 32732 25906
rect 32680 25842 32732 25848
rect 33428 25838 33456 26930
rect 33704 26382 33732 28086
rect 33784 26920 33836 26926
rect 33784 26862 33836 26868
rect 33980 26874 34008 34496
rect 35808 34478 35860 34484
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 36268 33992 36320 33998
rect 36268 33934 36320 33940
rect 36280 33522 36308 33934
rect 34704 33516 34756 33522
rect 34704 33458 34756 33464
rect 36268 33516 36320 33522
rect 36268 33458 36320 33464
rect 34716 32910 34744 33458
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34704 32904 34756 32910
rect 34704 32846 34756 32852
rect 36268 32904 36320 32910
rect 36268 32846 36320 32852
rect 34060 32768 34112 32774
rect 34060 32710 34112 32716
rect 34796 32768 34848 32774
rect 34796 32710 34848 32716
rect 34072 31890 34100 32710
rect 34704 32564 34756 32570
rect 34704 32506 34756 32512
rect 34152 32360 34204 32366
rect 34152 32302 34204 32308
rect 34164 31890 34192 32302
rect 34612 32020 34664 32026
rect 34612 31962 34664 31968
rect 34060 31884 34112 31890
rect 34060 31826 34112 31832
rect 34152 31884 34204 31890
rect 34152 31826 34204 31832
rect 34624 31346 34652 31962
rect 34716 31890 34744 32506
rect 34808 32434 34836 32710
rect 36280 32434 36308 32846
rect 34796 32428 34848 32434
rect 34796 32370 34848 32376
rect 36268 32428 36320 32434
rect 36268 32370 36320 32376
rect 36268 32224 36320 32230
rect 36268 32166 36320 32172
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 36280 31890 36308 32166
rect 34704 31884 34756 31890
rect 34704 31826 34756 31832
rect 36268 31884 36320 31890
rect 36268 31826 36320 31832
rect 36452 31748 36504 31754
rect 36452 31690 36504 31696
rect 36464 31482 36492 31690
rect 36452 31476 36504 31482
rect 36452 31418 36504 31424
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 36912 31340 36964 31346
rect 36912 31282 36964 31288
rect 34624 30734 34652 31282
rect 35440 31136 35492 31142
rect 35440 31078 35492 31084
rect 36084 31136 36136 31142
rect 36084 31078 36136 31084
rect 36452 31136 36504 31142
rect 36452 31078 36504 31084
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35452 30802 35480 31078
rect 35440 30796 35492 30802
rect 35440 30738 35492 30744
rect 34244 30728 34296 30734
rect 34244 30670 34296 30676
rect 34612 30728 34664 30734
rect 34612 30670 34664 30676
rect 35532 30728 35584 30734
rect 35532 30670 35584 30676
rect 34256 30190 34284 30670
rect 35256 30592 35308 30598
rect 35256 30534 35308 30540
rect 35268 30326 35296 30534
rect 35544 30394 35572 30670
rect 35532 30388 35584 30394
rect 35532 30330 35584 30336
rect 35256 30320 35308 30326
rect 35256 30262 35308 30268
rect 34244 30184 34296 30190
rect 34244 30126 34296 30132
rect 34256 29170 34284 30126
rect 34612 30048 34664 30054
rect 34612 29990 34664 29996
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 34244 29164 34296 29170
rect 34244 29106 34296 29112
rect 34060 28960 34112 28966
rect 34060 28902 34112 28908
rect 34152 28960 34204 28966
rect 34152 28902 34204 28908
rect 34072 28490 34100 28902
rect 34164 28762 34192 28902
rect 34152 28756 34204 28762
rect 34152 28698 34204 28704
rect 34532 28558 34560 29446
rect 34624 28762 34652 29990
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35544 29646 35572 30330
rect 36096 29714 36124 31078
rect 36464 30802 36492 31078
rect 36924 30938 36952 31282
rect 36912 30932 36964 30938
rect 36912 30874 36964 30880
rect 36452 30796 36504 30802
rect 36452 30738 36504 30744
rect 36544 30048 36596 30054
rect 36544 29990 36596 29996
rect 36084 29708 36136 29714
rect 36084 29650 36136 29656
rect 35532 29640 35584 29646
rect 35532 29582 35584 29588
rect 34704 29572 34756 29578
rect 34704 29514 34756 29520
rect 35348 29572 35400 29578
rect 35348 29514 35400 29520
rect 34612 28756 34664 28762
rect 34612 28698 34664 28704
rect 34520 28552 34572 28558
rect 34520 28494 34572 28500
rect 34060 28484 34112 28490
rect 34060 28426 34112 28432
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34428 27532 34480 27538
rect 34428 27474 34480 27480
rect 34336 27056 34388 27062
rect 34336 26998 34388 27004
rect 33692 26376 33744 26382
rect 33692 26318 33744 26324
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33416 25832 33468 25838
rect 33416 25774 33468 25780
rect 33612 25294 33640 25978
rect 32588 25288 32640 25294
rect 32588 25230 32640 25236
rect 33600 25288 33652 25294
rect 33600 25230 33652 25236
rect 32496 25220 32548 25226
rect 32496 25162 32548 25168
rect 31772 24670 31892 24698
rect 32404 24744 32456 24750
rect 32404 24686 32456 24692
rect 31392 24608 31444 24614
rect 31392 24550 31444 24556
rect 31404 24070 31432 24550
rect 31392 24064 31444 24070
rect 31392 24006 31444 24012
rect 31300 22976 31352 22982
rect 31300 22918 31352 22924
rect 31312 21690 31340 22918
rect 31300 21684 31352 21690
rect 31300 21626 31352 21632
rect 31484 20460 31536 20466
rect 31484 20402 31536 20408
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31298 20360 31354 20369
rect 31298 20295 31300 20304
rect 31352 20295 31354 20304
rect 31392 20324 31444 20330
rect 31300 20266 31352 20272
rect 31392 20266 31444 20272
rect 31208 18896 31260 18902
rect 31208 18838 31260 18844
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 31024 18692 31076 18698
rect 30944 18652 31024 18680
rect 30656 18352 30708 18358
rect 30656 18294 30708 18300
rect 30656 17808 30708 17814
rect 30656 17750 30708 17756
rect 30288 16788 30340 16794
rect 30288 16730 30340 16736
rect 30196 16720 30248 16726
rect 30196 16662 30248 16668
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30208 15570 30236 16662
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30288 16040 30340 16046
rect 30288 15982 30340 15988
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30300 15162 30328 15982
rect 30392 15502 30420 16458
rect 30472 16448 30524 16454
rect 30472 16390 30524 16396
rect 30484 15978 30512 16390
rect 30472 15972 30524 15978
rect 30472 15914 30524 15920
rect 30484 15502 30512 15914
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 30484 15178 30512 15438
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29828 15156 29880 15162
rect 29828 15098 29880 15104
rect 30288 15156 30340 15162
rect 30288 15098 30340 15104
rect 30392 15150 30512 15178
rect 29144 14980 29224 15008
rect 29092 14962 29144 14968
rect 29000 14816 29052 14822
rect 29000 14758 29052 14764
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28632 14000 28684 14006
rect 28632 13942 28684 13948
rect 28644 13870 28672 13942
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 27896 13524 27948 13530
rect 27896 13466 27948 13472
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27712 12640 27764 12646
rect 27712 12582 27764 12588
rect 27620 12164 27672 12170
rect 27620 12106 27672 12112
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27264 11014 27292 11154
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 26976 10736 27028 10742
rect 26976 10678 27028 10684
rect 27264 10674 27292 10950
rect 27632 10810 27660 12106
rect 27724 11694 27752 12582
rect 27712 11688 27764 11694
rect 27712 11630 27764 11636
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27816 10266 27844 11086
rect 27908 11014 27936 13466
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28644 12918 28672 13194
rect 28632 12912 28684 12918
rect 28632 12854 28684 12860
rect 28828 12442 28856 14214
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 29012 12238 29040 14758
rect 29380 13870 29408 15098
rect 30392 15042 30420 15150
rect 29552 15020 29604 15026
rect 29552 14962 29604 14968
rect 30300 15014 30420 15042
rect 29564 14482 29592 14962
rect 30300 14482 30328 15014
rect 30576 14822 30604 15302
rect 30564 14816 30616 14822
rect 30564 14758 30616 14764
rect 29552 14476 29604 14482
rect 29552 14418 29604 14424
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 30576 14074 30604 14758
rect 29552 14068 29604 14074
rect 29472 14028 29552 14056
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 29472 13394 29500 14028
rect 29552 14010 29604 14016
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 29920 13864 29972 13870
rect 29920 13806 29972 13812
rect 29552 13728 29604 13734
rect 29552 13670 29604 13676
rect 29276 13388 29328 13394
rect 29276 13330 29328 13336
rect 29460 13388 29512 13394
rect 29460 13330 29512 13336
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28632 11552 28684 11558
rect 28632 11494 28684 11500
rect 27896 11008 27948 11014
rect 27896 10950 27948 10956
rect 28172 10736 28224 10742
rect 28172 10678 28224 10684
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 27804 10260 27856 10266
rect 27804 10202 27856 10208
rect 27896 10260 27948 10266
rect 27896 10202 27948 10208
rect 27540 10130 27752 10146
rect 27528 10124 27752 10130
rect 27580 10118 27752 10124
rect 27528 10066 27580 10072
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 27172 9654 27568 9674
rect 27172 9648 27580 9654
rect 27172 9646 27528 9648
rect 27172 9586 27200 9646
rect 27528 9590 27580 9596
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 26516 9512 26568 9518
rect 26516 9454 26568 9460
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26292 8792 26372 8820
rect 26240 8774 26292 8780
rect 26344 8498 26372 8792
rect 26424 8832 26476 8838
rect 26424 8774 26476 8780
rect 26436 8566 26464 8774
rect 26424 8560 26476 8566
rect 26424 8502 26476 8508
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 26344 7954 26372 8434
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26436 8022 26464 8366
rect 26424 8016 26476 8022
rect 26424 7958 26476 7964
rect 26332 7948 26384 7954
rect 26332 7890 26384 7896
rect 26436 7546 26464 7958
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 25780 7404 25832 7410
rect 25780 7346 25832 7352
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 25688 5296 25740 5302
rect 25688 5238 25740 5244
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24504 4214 24532 4422
rect 24492 4208 24544 4214
rect 24492 4150 24544 4156
rect 24780 4146 24808 4626
rect 25700 4146 25728 5238
rect 25792 4486 25820 5646
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 25884 5302 25912 5510
rect 25872 5296 25924 5302
rect 25872 5238 25924 5244
rect 25976 4554 26004 5510
rect 26252 4554 26280 7142
rect 26344 7041 26372 7346
rect 26330 7032 26386 7041
rect 26330 6967 26386 6976
rect 26344 6798 26372 6967
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26528 6322 26556 9454
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26792 8832 26844 8838
rect 26792 8774 26844 8780
rect 26804 7818 26832 8774
rect 26896 8634 26924 8842
rect 26884 8628 26936 8634
rect 26884 8570 26936 8576
rect 26988 7886 27016 9318
rect 27172 7886 27200 9522
rect 27448 9110 27476 9522
rect 27436 9104 27488 9110
rect 27436 9046 27488 9052
rect 27436 8900 27488 8906
rect 27436 8842 27488 8848
rect 26976 7880 27028 7886
rect 27160 7880 27212 7886
rect 26976 7822 27028 7828
rect 27158 7848 27160 7857
rect 27212 7848 27214 7857
rect 26792 7812 26844 7818
rect 27158 7783 27214 7792
rect 27252 7812 27304 7818
rect 26792 7754 26844 7760
rect 27252 7754 27304 7760
rect 26804 7002 26832 7754
rect 27264 7546 27292 7754
rect 27448 7562 27476 8842
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27632 8498 27660 8774
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27632 8362 27660 8434
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27540 7886 27568 7958
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27632 7750 27660 8298
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27356 7534 27476 7562
rect 27356 7410 27384 7534
rect 27434 7440 27490 7449
rect 27068 7404 27120 7410
rect 27068 7346 27120 7352
rect 27344 7404 27396 7410
rect 27434 7375 27490 7384
rect 27344 7346 27396 7352
rect 26976 7200 27028 7206
rect 26976 7142 27028 7148
rect 26792 6996 26844 7002
rect 26792 6938 26844 6944
rect 26988 6798 27016 7142
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 27080 6458 27108 7346
rect 27448 7342 27476 7375
rect 27724 7342 27752 10118
rect 27908 10062 27936 10202
rect 28092 10062 28120 10610
rect 28184 10606 28212 10678
rect 28644 10674 28672 11494
rect 28632 10668 28684 10674
rect 28632 10610 28684 10616
rect 28172 10600 28224 10606
rect 28172 10542 28224 10548
rect 28184 10130 28212 10542
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 27896 10056 27948 10062
rect 27816 10016 27896 10044
rect 27816 8974 27844 10016
rect 27896 9998 27948 10004
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 27908 9518 27936 9862
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27988 8900 28040 8906
rect 27988 8842 28040 8848
rect 28000 8809 28028 8842
rect 28092 8838 28120 9998
rect 28276 9722 28304 9998
rect 28540 9988 28592 9994
rect 28540 9930 28592 9936
rect 28264 9716 28316 9722
rect 28264 9658 28316 9664
rect 28276 8974 28304 9658
rect 28552 9110 28580 9930
rect 28632 9512 28684 9518
rect 28736 9466 28764 11630
rect 29184 11280 29236 11286
rect 29184 11222 29236 11228
rect 29196 10810 29224 11222
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 29288 10742 29316 13330
rect 29564 12850 29592 13670
rect 29932 13530 29960 13806
rect 30668 13530 30696 17750
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 30760 16998 30788 17478
rect 30748 16992 30800 16998
rect 30748 16934 30800 16940
rect 30944 16590 30972 18652
rect 31024 18634 31076 18640
rect 31116 18624 31168 18630
rect 31116 18566 31168 18572
rect 31024 18420 31076 18426
rect 31024 18362 31076 18368
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 31036 16522 31064 18362
rect 31128 18086 31156 18566
rect 31116 18080 31168 18086
rect 31116 18022 31168 18028
rect 31116 17128 31168 17134
rect 31116 17070 31168 17076
rect 31024 16516 31076 16522
rect 31024 16458 31076 16464
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30760 16114 30788 16390
rect 31128 16250 31156 17070
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 30760 15116 30972 15144
rect 30760 14550 30788 15116
rect 30944 15076 30972 15116
rect 31220 15094 31248 15438
rect 31024 15088 31076 15094
rect 30944 15048 31024 15076
rect 31024 15030 31076 15036
rect 31208 15088 31260 15094
rect 31208 15030 31260 15036
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 31116 15020 31168 15026
rect 31116 14962 31168 14968
rect 30748 14544 30800 14550
rect 30748 14486 30800 14492
rect 29644 13524 29696 13530
rect 29644 13466 29696 13472
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 30656 13524 30708 13530
rect 30656 13466 30708 13472
rect 29552 12844 29604 12850
rect 29552 12786 29604 12792
rect 29656 12782 29684 13466
rect 30760 13258 30788 14486
rect 30852 14414 30880 14962
rect 31024 14816 31076 14822
rect 31024 14758 31076 14764
rect 30840 14408 30892 14414
rect 30892 14368 30972 14396
rect 30840 14350 30892 14356
rect 30748 13252 30800 13258
rect 30748 13194 30800 13200
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30286 12880 30342 12889
rect 29736 12844 29788 12850
rect 29736 12786 29788 12792
rect 29920 12844 29972 12850
rect 30286 12815 30342 12824
rect 29920 12786 29972 12792
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29460 12640 29512 12646
rect 29460 12582 29512 12588
rect 29368 12096 29420 12102
rect 29368 12038 29420 12044
rect 29380 11218 29408 12038
rect 29472 11830 29500 12582
rect 29748 12442 29776 12786
rect 29932 12442 29960 12786
rect 30300 12714 30328 12815
rect 30288 12708 30340 12714
rect 30288 12650 30340 12656
rect 30380 12708 30432 12714
rect 30380 12650 30432 12656
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29920 12436 29972 12442
rect 29920 12378 29972 12384
rect 30392 12238 30420 12650
rect 30484 12238 30512 13126
rect 30944 12850 30972 14368
rect 31036 14074 31064 14758
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 31036 13394 31064 14010
rect 31128 14006 31156 14962
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 31220 14074 31248 14350
rect 31208 14068 31260 14074
rect 31208 14010 31260 14016
rect 31116 14000 31168 14006
rect 31116 13942 31168 13948
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 31116 13864 31168 13870
rect 31116 13806 31168 13812
rect 31024 13388 31076 13394
rect 31024 13330 31076 13336
rect 31024 13252 31076 13258
rect 31024 13194 31076 13200
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 30944 12238 30972 12786
rect 31036 12238 31064 13194
rect 31128 12782 31156 13806
rect 31220 13326 31248 13874
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31220 12850 31248 13262
rect 31312 12918 31340 20266
rect 31404 20058 31432 20266
rect 31392 20052 31444 20058
rect 31392 19994 31444 20000
rect 31496 19825 31524 20402
rect 31482 19816 31538 19825
rect 31680 19786 31708 20402
rect 31482 19751 31538 19760
rect 31668 19780 31720 19786
rect 31668 19722 31720 19728
rect 31484 19304 31536 19310
rect 31484 19246 31536 19252
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 31392 18964 31444 18970
rect 31392 18906 31444 18912
rect 31404 17542 31432 18906
rect 31496 18290 31524 19246
rect 31588 18970 31616 19246
rect 31576 18964 31628 18970
rect 31576 18906 31628 18912
rect 31680 18426 31708 19722
rect 31668 18420 31720 18426
rect 31668 18362 31720 18368
rect 31484 18284 31536 18290
rect 31484 18226 31536 18232
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 31496 16590 31524 18226
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 31680 17134 31708 18158
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31484 16584 31536 16590
rect 31484 16526 31536 16532
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31404 13190 31432 16050
rect 31680 15910 31708 17070
rect 31668 15904 31720 15910
rect 31668 15846 31720 15852
rect 31680 15570 31708 15846
rect 31668 15564 31720 15570
rect 31668 15506 31720 15512
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 31496 15162 31524 15438
rect 31484 15156 31536 15162
rect 31484 15098 31536 15104
rect 31680 15026 31708 15506
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31484 14952 31536 14958
rect 31484 14894 31536 14900
rect 31496 14482 31524 14894
rect 31772 14550 31800 24670
rect 32036 24608 32088 24614
rect 32036 24550 32088 24556
rect 31944 24200 31996 24206
rect 31944 24142 31996 24148
rect 31956 23594 31984 24142
rect 31944 23588 31996 23594
rect 31944 23530 31996 23536
rect 32048 23186 32076 24550
rect 32508 24410 32536 25162
rect 33508 24812 33560 24818
rect 33508 24754 33560 24760
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 32496 24404 32548 24410
rect 32496 24346 32548 24352
rect 32968 24342 32996 24686
rect 33520 24410 33548 24754
rect 33796 24750 33824 26862
rect 33876 26852 33928 26858
rect 33980 26846 34192 26874
rect 33876 26794 33928 26800
rect 33888 26314 33916 26794
rect 34060 26784 34112 26790
rect 34060 26726 34112 26732
rect 34072 26382 34100 26726
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 34060 26376 34112 26382
rect 34060 26318 34112 26324
rect 33876 26308 33928 26314
rect 33876 26250 33928 26256
rect 33980 26042 34008 26318
rect 33968 26036 34020 26042
rect 33968 25978 34020 25984
rect 34072 25226 34100 26318
rect 34060 25220 34112 25226
rect 34060 25162 34112 25168
rect 34164 25106 34192 26846
rect 34348 25906 34376 26998
rect 34440 26586 34468 27474
rect 34532 27062 34560 27950
rect 34612 27872 34664 27878
rect 34612 27814 34664 27820
rect 34624 27606 34652 27814
rect 34612 27600 34664 27606
rect 34612 27542 34664 27548
rect 34716 27334 34744 29514
rect 35360 29102 35388 29514
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 35348 29096 35400 29102
rect 35348 29038 35400 29044
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35360 28626 35388 29038
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 35348 28620 35400 28626
rect 35348 28562 35400 28568
rect 34808 28422 34836 28562
rect 34980 28552 35032 28558
rect 34980 28494 35032 28500
rect 34796 28416 34848 28422
rect 34796 28358 34848 28364
rect 34992 28218 35020 28494
rect 35716 28416 35768 28422
rect 35716 28358 35768 28364
rect 34888 28212 34940 28218
rect 34808 28172 34888 28200
rect 34704 27328 34756 27334
rect 34704 27270 34756 27276
rect 34520 27056 34572 27062
rect 34520 26998 34572 27004
rect 34716 26994 34744 27270
rect 34808 27130 34836 28172
rect 34888 28154 34940 28160
rect 34980 28212 35032 28218
rect 34980 28154 35032 28160
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35532 27396 35584 27402
rect 35532 27338 35584 27344
rect 34796 27124 34848 27130
rect 34796 27066 34848 27072
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34428 26580 34480 26586
rect 34428 26522 34480 26528
rect 34612 26512 34664 26518
rect 34612 26454 34664 26460
rect 34624 25974 34652 26454
rect 34808 26450 34836 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34796 26444 34848 26450
rect 34796 26386 34848 26392
rect 35452 26382 35480 26930
rect 35544 26382 35572 27338
rect 35624 26920 35676 26926
rect 35624 26862 35676 26868
rect 35440 26376 35492 26382
rect 35440 26318 35492 26324
rect 35532 26376 35584 26382
rect 35532 26318 35584 26324
rect 35452 26042 35480 26318
rect 35636 26314 35664 26862
rect 35624 26308 35676 26314
rect 35624 26250 35676 26256
rect 35440 26036 35492 26042
rect 35440 25978 35492 25984
rect 34612 25968 34664 25974
rect 34612 25910 34664 25916
rect 35348 25968 35400 25974
rect 35348 25910 35400 25916
rect 34336 25900 34388 25906
rect 34336 25842 34388 25848
rect 34072 25078 34192 25106
rect 33784 24744 33836 24750
rect 33784 24686 33836 24692
rect 33508 24404 33560 24410
rect 33508 24346 33560 24352
rect 32956 24336 33008 24342
rect 32956 24278 33008 24284
rect 33508 24268 33560 24274
rect 33508 24210 33560 24216
rect 32772 24132 32824 24138
rect 32772 24074 32824 24080
rect 32784 23866 32812 24074
rect 32772 23860 32824 23866
rect 32772 23802 32824 23808
rect 33520 23730 33548 24210
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 33692 23656 33744 23662
rect 33692 23598 33744 23604
rect 32036 23180 32088 23186
rect 32036 23122 32088 23128
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31864 21622 31892 22986
rect 31944 22500 31996 22506
rect 31944 22442 31996 22448
rect 31852 21616 31904 21622
rect 31852 21558 31904 21564
rect 31956 20874 31984 22442
rect 32048 21010 32076 23122
rect 33416 23112 33468 23118
rect 33416 23054 33468 23060
rect 32312 23044 32364 23050
rect 32312 22986 32364 22992
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32140 21962 32168 22374
rect 32128 21956 32180 21962
rect 32128 21898 32180 21904
rect 32220 21888 32272 21894
rect 32220 21830 32272 21836
rect 32232 21434 32260 21830
rect 32140 21406 32260 21434
rect 32036 21004 32088 21010
rect 32036 20946 32088 20952
rect 31944 20868 31996 20874
rect 31944 20810 31996 20816
rect 32140 20398 32168 21406
rect 32220 21344 32272 21350
rect 32220 21286 32272 21292
rect 32128 20392 32180 20398
rect 32128 20334 32180 20340
rect 32232 19854 32260 21286
rect 32324 20058 32352 22986
rect 33048 22976 33100 22982
rect 33048 22918 33100 22924
rect 33060 22234 33088 22918
rect 33428 22778 33456 23054
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 33060 22094 33088 22170
rect 32968 22066 33088 22094
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32312 20052 32364 20058
rect 32312 19994 32364 20000
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32048 18873 32076 19790
rect 32416 19530 32444 21490
rect 32588 20528 32640 20534
rect 32588 20470 32640 20476
rect 32496 19984 32548 19990
rect 32496 19926 32548 19932
rect 32324 19502 32444 19530
rect 32324 19310 32352 19502
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 32324 19174 32352 19246
rect 32508 19174 32536 19926
rect 32220 19168 32272 19174
rect 32220 19110 32272 19116
rect 32312 19168 32364 19174
rect 32312 19110 32364 19116
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32034 18864 32090 18873
rect 32034 18799 32090 18808
rect 32232 18766 32260 19110
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32496 18692 32548 18698
rect 32496 18634 32548 18640
rect 32404 18624 32456 18630
rect 32404 18566 32456 18572
rect 32416 18154 32444 18566
rect 32404 18148 32456 18154
rect 32404 18090 32456 18096
rect 32508 17542 32536 18634
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32496 17536 32548 17542
rect 32496 17478 32548 17484
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31944 16720 31996 16726
rect 31944 16662 31996 16668
rect 31956 16561 31984 16662
rect 31942 16552 31998 16561
rect 31942 16487 31998 16496
rect 31760 14544 31812 14550
rect 31760 14486 31812 14492
rect 31484 14476 31536 14482
rect 31484 14418 31536 14424
rect 31496 13818 31524 14418
rect 32048 14414 32076 17274
rect 32416 17066 32444 17478
rect 32404 17060 32456 17066
rect 32404 17002 32456 17008
rect 32128 16992 32180 16998
rect 32128 16934 32180 16940
rect 32140 16794 32168 16934
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 32220 16516 32272 16522
rect 32220 16458 32272 16464
rect 32232 14958 32260 16458
rect 32508 16454 32536 17478
rect 32496 16448 32548 16454
rect 32496 16390 32548 16396
rect 32600 16046 32628 20470
rect 32968 19854 32996 22066
rect 33232 21888 33284 21894
rect 33232 21830 33284 21836
rect 33244 21554 33272 21830
rect 33232 21548 33284 21554
rect 33232 21490 33284 21496
rect 33416 21548 33468 21554
rect 33416 21490 33468 21496
rect 33048 21480 33100 21486
rect 33048 21422 33100 21428
rect 33060 21010 33088 21422
rect 33428 21146 33456 21490
rect 33704 21146 33732 23598
rect 33876 22568 33928 22574
rect 33876 22510 33928 22516
rect 33784 22500 33836 22506
rect 33784 22442 33836 22448
rect 33796 22234 33824 22442
rect 33784 22228 33836 22234
rect 33784 22170 33836 22176
rect 33796 21146 33824 22170
rect 33416 21140 33468 21146
rect 33416 21082 33468 21088
rect 33692 21140 33744 21146
rect 33692 21082 33744 21088
rect 33784 21140 33836 21146
rect 33784 21082 33836 21088
rect 33048 21004 33100 21010
rect 33048 20946 33100 20952
rect 33140 20936 33192 20942
rect 33140 20878 33192 20884
rect 32956 19848 33008 19854
rect 32956 19790 33008 19796
rect 32968 19446 32996 19790
rect 32956 19440 33008 19446
rect 32956 19382 33008 19388
rect 32968 18426 32996 19382
rect 33152 19378 33180 20878
rect 33416 20868 33468 20874
rect 33416 20810 33468 20816
rect 33428 20602 33456 20810
rect 33416 20596 33468 20602
rect 33416 20538 33468 20544
rect 33888 20466 33916 22510
rect 34072 22094 34100 25078
rect 34348 24818 34376 25842
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35360 25498 35388 25910
rect 35636 25838 35664 26250
rect 35624 25832 35676 25838
rect 35624 25774 35676 25780
rect 35348 25492 35400 25498
rect 35348 25434 35400 25440
rect 35728 25362 35756 28358
rect 35912 28082 35940 29446
rect 36556 29238 36584 29990
rect 36544 29232 36596 29238
rect 36544 29174 36596 29180
rect 35900 28076 35952 28082
rect 35900 28018 35952 28024
rect 36268 27464 36320 27470
rect 36268 27406 36320 27412
rect 36280 26897 36308 27406
rect 36266 26888 36322 26897
rect 36266 26823 36322 26832
rect 35808 26376 35860 26382
rect 35808 26318 35860 26324
rect 36268 26376 36320 26382
rect 36268 26318 36320 26324
rect 35716 25356 35768 25362
rect 35716 25298 35768 25304
rect 35348 25288 35400 25294
rect 35348 25230 35400 25236
rect 34612 25152 34664 25158
rect 34612 25094 34664 25100
rect 34336 24812 34388 24818
rect 34336 24754 34388 24760
rect 34348 24682 34376 24754
rect 34624 24750 34652 25094
rect 34612 24744 34664 24750
rect 34612 24686 34664 24692
rect 34336 24676 34388 24682
rect 34336 24618 34388 24624
rect 34348 23798 34376 24618
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34704 24336 34756 24342
rect 34704 24278 34756 24284
rect 34716 24206 34744 24278
rect 35360 24206 35388 25230
rect 35716 24812 35768 24818
rect 35716 24754 35768 24760
rect 35728 24410 35756 24754
rect 35820 24750 35848 26318
rect 36280 25362 36308 26318
rect 36452 25696 36504 25702
rect 36452 25638 36504 25644
rect 36464 25362 36492 25638
rect 36268 25356 36320 25362
rect 36268 25298 36320 25304
rect 36452 25356 36504 25362
rect 36452 25298 36504 25304
rect 35808 24744 35860 24750
rect 35808 24686 35860 24692
rect 36268 24608 36320 24614
rect 36268 24550 36320 24556
rect 35716 24404 35768 24410
rect 35716 24346 35768 24352
rect 36280 24274 36308 24550
rect 36268 24268 36320 24274
rect 36268 24210 36320 24216
rect 34612 24200 34664 24206
rect 34612 24142 34664 24148
rect 34704 24200 34756 24206
rect 34704 24142 34756 24148
rect 35348 24200 35400 24206
rect 35348 24142 35400 24148
rect 35440 24200 35492 24206
rect 35440 24142 35492 24148
rect 34428 24132 34480 24138
rect 34428 24074 34480 24080
rect 34520 24132 34572 24138
rect 34520 24074 34572 24080
rect 34336 23792 34388 23798
rect 34336 23734 34388 23740
rect 34336 23656 34388 23662
rect 34440 23610 34468 24074
rect 34532 23866 34560 24074
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34388 23604 34468 23610
rect 34336 23598 34468 23604
rect 34348 23582 34468 23598
rect 34520 23316 34572 23322
rect 34520 23258 34572 23264
rect 34072 22066 34284 22094
rect 33968 21888 34020 21894
rect 33968 21830 34020 21836
rect 34060 21888 34112 21894
rect 34060 21830 34112 21836
rect 33980 20534 34008 21830
rect 34072 21554 34100 21830
rect 34060 21548 34112 21554
rect 34060 21490 34112 21496
rect 33968 20528 34020 20534
rect 33968 20470 34020 20476
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33324 19712 33376 19718
rect 33324 19654 33376 19660
rect 33336 19514 33364 19654
rect 33324 19508 33376 19514
rect 33324 19450 33376 19456
rect 33428 19378 33456 19790
rect 33508 19712 33560 19718
rect 33508 19654 33560 19660
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33416 19372 33468 19378
rect 33416 19314 33468 19320
rect 33232 19168 33284 19174
rect 33232 19110 33284 19116
rect 33048 18760 33100 18766
rect 33048 18702 33100 18708
rect 32956 18420 33008 18426
rect 32956 18362 33008 18368
rect 33060 18290 33088 18702
rect 33244 18698 33272 19110
rect 33232 18692 33284 18698
rect 33232 18634 33284 18640
rect 33324 18692 33376 18698
rect 33324 18634 33376 18640
rect 33140 18624 33192 18630
rect 33140 18566 33192 18572
rect 32864 18284 32916 18290
rect 32864 18226 32916 18232
rect 33048 18284 33100 18290
rect 33048 18226 33100 18232
rect 32876 18170 32904 18226
rect 32680 18148 32732 18154
rect 32876 18142 32996 18170
rect 32680 18090 32732 18096
rect 32692 17270 32720 18090
rect 32968 18086 32996 18142
rect 32956 18080 33008 18086
rect 32956 18022 33008 18028
rect 32864 17876 32916 17882
rect 32864 17818 32916 17824
rect 32772 17808 32824 17814
rect 32772 17750 32824 17756
rect 32680 17264 32732 17270
rect 32680 17206 32732 17212
rect 32784 16590 32812 17750
rect 32876 17338 32904 17818
rect 32968 17610 32996 18022
rect 33060 17882 33088 18226
rect 33048 17876 33100 17882
rect 33048 17818 33100 17824
rect 32956 17604 33008 17610
rect 32956 17546 33008 17552
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 32968 16998 32996 17546
rect 33152 17338 33180 18566
rect 33230 18048 33286 18057
rect 33230 17983 33286 17992
rect 33244 17678 33272 17983
rect 33232 17672 33284 17678
rect 33232 17614 33284 17620
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 33048 17264 33100 17270
rect 33048 17206 33100 17212
rect 32956 16992 33008 16998
rect 32956 16934 33008 16940
rect 33060 16590 33088 17206
rect 32772 16584 32824 16590
rect 32772 16526 32824 16532
rect 33048 16584 33100 16590
rect 33048 16526 33100 16532
rect 33140 16176 33192 16182
rect 33140 16118 33192 16124
rect 32956 16108 33008 16114
rect 32956 16050 33008 16056
rect 32588 16040 32640 16046
rect 32588 15982 32640 15988
rect 32312 15632 32364 15638
rect 32364 15580 32444 15586
rect 32312 15574 32444 15580
rect 32324 15558 32444 15574
rect 32416 15162 32444 15558
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 32220 14952 32272 14958
rect 32220 14894 32272 14900
rect 32036 14408 32088 14414
rect 32036 14350 32088 14356
rect 31576 14272 31628 14278
rect 31576 14214 31628 14220
rect 31588 14006 31616 14214
rect 31576 14000 31628 14006
rect 31576 13942 31628 13948
rect 32048 13938 32076 14350
rect 32232 14346 32260 14894
rect 32416 14822 32444 15098
rect 32496 15088 32548 15094
rect 32496 15030 32548 15036
rect 32312 14816 32364 14822
rect 32312 14758 32364 14764
rect 32404 14816 32456 14822
rect 32404 14758 32456 14764
rect 32324 14618 32352 14758
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32220 14340 32272 14346
rect 32220 14282 32272 14288
rect 32036 13932 32088 13938
rect 32036 13874 32088 13880
rect 31576 13864 31628 13870
rect 31496 13812 31576 13818
rect 31496 13806 31628 13812
rect 31496 13790 31616 13806
rect 31392 13184 31444 13190
rect 31392 13126 31444 13132
rect 31300 12912 31352 12918
rect 31300 12854 31352 12860
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31116 12776 31168 12782
rect 31116 12718 31168 12724
rect 30380 12232 30432 12238
rect 30472 12232 30524 12238
rect 30380 12174 30432 12180
rect 30470 12200 30472 12209
rect 30932 12232 30984 12238
rect 30524 12200 30526 12209
rect 30932 12174 30984 12180
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 30470 12135 30526 12144
rect 30748 12164 30800 12170
rect 30484 12109 30512 12135
rect 30748 12106 30800 12112
rect 30760 11898 30788 12106
rect 30472 11892 30524 11898
rect 30472 11834 30524 11840
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 29460 11824 29512 11830
rect 29460 11766 29512 11772
rect 29920 11824 29972 11830
rect 29920 11766 29972 11772
rect 29932 11354 29960 11766
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 29368 11212 29420 11218
rect 29368 11154 29420 11160
rect 29276 10736 29328 10742
rect 29276 10678 29328 10684
rect 29380 10470 29408 11154
rect 30380 11144 30432 11150
rect 30380 11086 30432 11092
rect 30392 10810 30420 11086
rect 30380 10804 30432 10810
rect 30380 10746 30432 10752
rect 29828 10736 29880 10742
rect 29828 10678 29880 10684
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 29000 10192 29052 10198
rect 29000 10134 29052 10140
rect 29012 9994 29040 10134
rect 29840 10062 29868 10678
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 30208 10266 30236 10542
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 29644 10056 29696 10062
rect 29644 9998 29696 10004
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 28684 9460 28764 9466
rect 28632 9454 28764 9460
rect 28644 9438 28764 9454
rect 28540 9104 28592 9110
rect 28540 9046 28592 9052
rect 28264 8968 28316 8974
rect 28264 8910 28316 8916
rect 28080 8832 28132 8838
rect 27986 8800 28042 8809
rect 28080 8774 28132 8780
rect 27986 8735 28042 8744
rect 27804 8628 27856 8634
rect 27804 8570 27856 8576
rect 27816 8430 27844 8570
rect 27804 8424 27856 8430
rect 27804 8366 27856 8372
rect 27804 8016 27856 8022
rect 27802 7984 27804 7993
rect 27856 7984 27858 7993
rect 27802 7919 27858 7928
rect 28276 7886 28304 8910
rect 28736 8430 28764 9438
rect 29656 8974 29684 9998
rect 30208 9722 30236 10202
rect 30392 10062 30420 10746
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 30012 9580 30064 9586
rect 30012 9522 30064 9528
rect 30024 9178 30052 9522
rect 30012 9172 30064 9178
rect 30012 9114 30064 9120
rect 30392 8974 30420 9862
rect 30484 9654 30512 11834
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30852 10742 30880 11494
rect 30944 11354 30972 12174
rect 31128 12102 31156 12718
rect 31220 12170 31248 12786
rect 31208 12164 31260 12170
rect 31208 12106 31260 12112
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 31220 11626 31248 12106
rect 31208 11620 31260 11626
rect 31208 11562 31260 11568
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 30932 11076 30984 11082
rect 30932 11018 30984 11024
rect 30840 10736 30892 10742
rect 30840 10678 30892 10684
rect 30944 10266 30972 11018
rect 31024 11008 31076 11014
rect 31024 10950 31076 10956
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 31036 9994 31064 10950
rect 31404 10742 31432 13126
rect 31588 11898 31616 13790
rect 32048 12918 32076 13874
rect 32508 13394 32536 15030
rect 32600 13734 32628 15982
rect 32968 15910 32996 16050
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 32968 13938 32996 15846
rect 33152 15706 33180 16118
rect 33140 15700 33192 15706
rect 33140 15642 33192 15648
rect 33244 13938 33272 17614
rect 33336 16522 33364 18634
rect 33520 18426 33548 19654
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33508 18420 33560 18426
rect 33508 18362 33560 18368
rect 33704 17678 33732 18566
rect 33692 17672 33744 17678
rect 33692 17614 33744 17620
rect 33600 17264 33652 17270
rect 33600 17206 33652 17212
rect 33324 16516 33376 16522
rect 33612 16504 33640 17206
rect 33704 16998 33732 17614
rect 33692 16992 33744 16998
rect 33692 16934 33744 16940
rect 33692 16516 33744 16522
rect 33612 16476 33692 16504
rect 33324 16458 33376 16464
rect 33692 16458 33744 16464
rect 33324 15904 33376 15910
rect 33324 15846 33376 15852
rect 33336 15094 33364 15846
rect 33324 15088 33376 15094
rect 33324 15030 33376 15036
rect 33600 14272 33652 14278
rect 33600 14214 33652 14220
rect 32956 13932 33008 13938
rect 32956 13874 33008 13880
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 32588 13728 32640 13734
rect 32588 13670 32640 13676
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32036 12912 32088 12918
rect 32404 12912 32456 12918
rect 32036 12854 32088 12860
rect 32402 12880 32404 12889
rect 32456 12880 32458 12889
rect 31852 12640 31904 12646
rect 31852 12582 31904 12588
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 31576 11892 31628 11898
rect 31576 11834 31628 11840
rect 31668 11688 31720 11694
rect 31668 11630 31720 11636
rect 31576 11552 31628 11558
rect 31576 11494 31628 11500
rect 31588 11082 31616 11494
rect 31680 11218 31708 11630
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31576 11076 31628 11082
rect 31576 11018 31628 11024
rect 31680 10810 31708 11154
rect 31668 10804 31720 10810
rect 31668 10746 31720 10752
rect 31392 10736 31444 10742
rect 31392 10678 31444 10684
rect 31668 10600 31720 10606
rect 31668 10542 31720 10548
rect 31680 10266 31708 10542
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31772 10062 31800 12038
rect 31864 11762 31892 12582
rect 32048 11830 32076 12854
rect 32402 12815 32458 12824
rect 32404 12776 32456 12782
rect 32404 12718 32456 12724
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32324 12442 32352 12582
rect 32312 12436 32364 12442
rect 32312 12378 32364 12384
rect 32416 12306 32444 12718
rect 32508 12714 32536 13330
rect 33612 12850 33640 14214
rect 33704 12918 33732 16458
rect 33796 14822 33824 19654
rect 33888 17814 33916 20402
rect 33980 19514 34008 20470
rect 33968 19508 34020 19514
rect 33968 19450 34020 19456
rect 33876 17808 33928 17814
rect 33876 17750 33928 17756
rect 33876 16788 33928 16794
rect 33876 16730 33928 16736
rect 33888 16182 33916 16730
rect 33876 16176 33928 16182
rect 33876 16118 33928 16124
rect 34060 16108 34112 16114
rect 34060 16050 34112 16056
rect 34072 15502 34100 16050
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 33784 14816 33836 14822
rect 33784 14758 33836 14764
rect 33876 14612 33928 14618
rect 33876 14554 33928 14560
rect 33888 13870 33916 14554
rect 34152 14408 34204 14414
rect 34152 14350 34204 14356
rect 33968 14340 34020 14346
rect 33968 14282 34020 14288
rect 33876 13864 33928 13870
rect 33876 13806 33928 13812
rect 33888 13462 33916 13806
rect 33876 13456 33928 13462
rect 33876 13398 33928 13404
rect 33980 13326 34008 14282
rect 34164 13938 34192 14350
rect 34152 13932 34204 13938
rect 34152 13874 34204 13880
rect 34152 13524 34204 13530
rect 34152 13466 34204 13472
rect 34060 13456 34112 13462
rect 34060 13398 34112 13404
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 33968 13320 34020 13326
rect 33968 13262 34020 13268
rect 33692 12912 33744 12918
rect 33692 12854 33744 12860
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 32496 12708 32548 12714
rect 32496 12650 32548 12656
rect 33612 12442 33640 12786
rect 33888 12782 33916 13262
rect 33876 12776 33928 12782
rect 33876 12718 33928 12724
rect 33600 12436 33652 12442
rect 33600 12378 33652 12384
rect 32494 12336 32550 12345
rect 32404 12300 32456 12306
rect 32494 12271 32550 12280
rect 32404 12242 32456 12248
rect 32416 12170 32444 12242
rect 32404 12164 32456 12170
rect 32404 12106 32456 12112
rect 32128 12096 32180 12102
rect 32128 12038 32180 12044
rect 32140 11898 32168 12038
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 32508 11830 32536 12271
rect 32680 12096 32732 12102
rect 32680 12038 32732 12044
rect 32036 11824 32088 11830
rect 32036 11766 32088 11772
rect 32496 11824 32548 11830
rect 32496 11766 32548 11772
rect 31852 11756 31904 11762
rect 31852 11698 31904 11704
rect 32692 11218 32720 12038
rect 32956 11756 33008 11762
rect 32956 11698 33008 11704
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 32128 10532 32180 10538
rect 32128 10474 32180 10480
rect 32140 10266 32168 10474
rect 32128 10260 32180 10266
rect 32128 10202 32180 10208
rect 32968 10062 32996 11698
rect 33416 11552 33468 11558
rect 33416 11494 33468 11500
rect 33428 10742 33456 11494
rect 33888 10810 33916 12718
rect 33980 12646 34008 13262
rect 34072 12986 34100 13398
rect 34164 13190 34192 13466
rect 34152 13184 34204 13190
rect 34152 13126 34204 13132
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 33968 12640 34020 12646
rect 33968 12582 34020 12588
rect 34164 12238 34192 13126
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 34164 11354 34192 12174
rect 34152 11348 34204 11354
rect 34152 11290 34204 11296
rect 33876 10804 33928 10810
rect 33876 10746 33928 10752
rect 33416 10736 33468 10742
rect 33416 10678 33468 10684
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 32956 10056 33008 10062
rect 32956 9998 33008 10004
rect 31024 9988 31076 9994
rect 31024 9930 31076 9936
rect 30472 9648 30524 9654
rect 30472 9590 30524 9596
rect 31036 9586 31064 9930
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 29656 8634 29684 8910
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 28724 8424 28776 8430
rect 28776 8372 28856 8378
rect 28724 8366 28856 8372
rect 28736 8350 28856 8366
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 27896 7812 27948 7818
rect 27896 7754 27948 7760
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 27816 7478 27844 7754
rect 27804 7472 27856 7478
rect 27804 7414 27856 7420
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27712 7336 27764 7342
rect 27712 7278 27764 7284
rect 27908 7002 27936 7754
rect 28460 7546 28488 7754
rect 28448 7540 28500 7546
rect 28448 7482 28500 7488
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 27068 6452 27120 6458
rect 27068 6394 27120 6400
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 27816 5914 27844 6326
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 28276 5166 28304 7278
rect 28540 6656 28592 6662
rect 28540 6598 28592 6604
rect 28552 6390 28580 6598
rect 28540 6384 28592 6390
rect 28540 6326 28592 6332
rect 28828 6322 28856 8350
rect 30208 7886 30236 8910
rect 30392 7886 30420 8910
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 30944 8090 30972 8502
rect 30932 8084 30984 8090
rect 30932 8026 30984 8032
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 30380 7880 30432 7886
rect 30380 7822 30432 7828
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 29012 6866 29040 7142
rect 29656 6866 29684 7346
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 29644 6860 29696 6866
rect 29644 6802 29696 6808
rect 30392 6798 30420 7822
rect 34256 6914 34284 22066
rect 34532 21690 34560 23258
rect 34624 22642 34652 24142
rect 34888 24064 34940 24070
rect 34888 24006 34940 24012
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 34900 23866 34928 24006
rect 34888 23860 34940 23866
rect 34888 23802 34940 23808
rect 35360 23730 35388 24006
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35452 23322 35480 24142
rect 35532 24064 35584 24070
rect 35532 24006 35584 24012
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 34704 22432 34756 22438
rect 34704 22374 34756 22380
rect 34520 21684 34572 21690
rect 34520 21626 34572 21632
rect 34716 21622 34744 22374
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35440 22160 35492 22166
rect 35440 22102 35492 22108
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34704 21616 34756 21622
rect 34704 21558 34756 21564
rect 34520 21412 34572 21418
rect 34520 21354 34572 21360
rect 34336 20460 34388 20466
rect 34336 20402 34388 20408
rect 34348 18970 34376 20402
rect 34532 20380 34560 21354
rect 34612 21344 34664 21350
rect 34612 21286 34664 21292
rect 34624 20534 34652 21286
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 34612 20528 34664 20534
rect 34612 20470 34664 20476
rect 34532 20352 34652 20380
rect 34428 20256 34480 20262
rect 34428 20198 34480 20204
rect 34520 20256 34572 20262
rect 34520 20198 34572 20204
rect 34440 19922 34468 20198
rect 34428 19916 34480 19922
rect 34428 19858 34480 19864
rect 34532 19446 34560 20198
rect 34520 19440 34572 19446
rect 34520 19382 34572 19388
rect 34520 19304 34572 19310
rect 34520 19246 34572 19252
rect 34428 19168 34480 19174
rect 34428 19110 34480 19116
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 34440 18698 34468 19110
rect 34532 18737 34560 19246
rect 34624 18986 34652 20352
rect 34716 19854 34744 20742
rect 34704 19848 34756 19854
rect 34704 19790 34756 19796
rect 34624 18958 34744 18986
rect 34518 18728 34574 18737
rect 34428 18692 34480 18698
rect 34518 18663 34574 18672
rect 34428 18634 34480 18640
rect 34520 18216 34572 18222
rect 34520 18158 34572 18164
rect 34612 18216 34664 18222
rect 34612 18158 34664 18164
rect 34532 17882 34560 18158
rect 34520 17876 34572 17882
rect 34520 17818 34572 17824
rect 34624 17338 34652 18158
rect 34612 17332 34664 17338
rect 34612 17274 34664 17280
rect 34716 16794 34744 18958
rect 34808 18766 34836 21966
rect 35348 21956 35400 21962
rect 35348 21898 35400 21904
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35360 20874 35388 21898
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 35360 20330 35388 20810
rect 35452 20516 35480 22102
rect 35544 20584 35572 24006
rect 36084 23588 36136 23594
rect 36084 23530 36136 23536
rect 35716 23520 35768 23526
rect 35716 23462 35768 23468
rect 35728 22234 35756 23462
rect 35992 23112 36044 23118
rect 35992 23054 36044 23060
rect 36004 22545 36032 23054
rect 35990 22536 36046 22545
rect 35990 22471 36046 22480
rect 36004 22234 36032 22471
rect 35716 22228 35768 22234
rect 35716 22170 35768 22176
rect 35992 22228 36044 22234
rect 35992 22170 36044 22176
rect 35728 21078 35756 22170
rect 35900 22092 35952 22098
rect 35900 22034 35952 22040
rect 35808 21684 35860 21690
rect 35808 21626 35860 21632
rect 35716 21072 35768 21078
rect 35716 21014 35768 21020
rect 35820 20618 35848 21626
rect 35912 20806 35940 22034
rect 36096 21622 36124 23530
rect 36360 23520 36412 23526
rect 36360 23462 36412 23468
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36372 23186 36400 23462
rect 36360 23180 36412 23186
rect 36360 23122 36412 23128
rect 36176 22976 36228 22982
rect 36176 22918 36228 22924
rect 36084 21616 36136 21622
rect 36084 21558 36136 21564
rect 35900 20800 35952 20806
rect 35900 20742 35952 20748
rect 35820 20590 35940 20618
rect 35544 20556 35756 20584
rect 35452 20488 35664 20516
rect 35348 20324 35400 20330
rect 35400 20284 35480 20312
rect 35348 20266 35400 20272
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35452 19854 35480 20284
rect 34980 19848 35032 19854
rect 34980 19790 35032 19796
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 34888 19712 34940 19718
rect 34888 19654 34940 19660
rect 34900 19310 34928 19654
rect 34888 19304 34940 19310
rect 34992 19281 35020 19790
rect 35532 19780 35584 19786
rect 35532 19722 35584 19728
rect 35348 19304 35400 19310
rect 34888 19246 34940 19252
rect 34978 19272 35034 19281
rect 35348 19246 35400 19252
rect 34978 19207 35034 19216
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34796 18760 34848 18766
rect 34796 18702 34848 18708
rect 34886 18728 34942 18737
rect 34886 18663 34942 18672
rect 34900 18630 34928 18663
rect 34796 18624 34848 18630
rect 34796 18566 34848 18572
rect 34888 18624 34940 18630
rect 34888 18566 34940 18572
rect 34808 18426 34836 18566
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 35360 17882 35388 19246
rect 35440 19168 35492 19174
rect 35438 19136 35440 19145
rect 35492 19136 35494 19145
rect 35438 19071 35494 19080
rect 35544 18986 35572 19722
rect 35452 18958 35572 18986
rect 35452 18630 35480 18958
rect 35532 18896 35584 18902
rect 35636 18850 35664 20488
rect 35728 20482 35756 20556
rect 35912 20516 35940 20590
rect 35912 20488 36032 20516
rect 35728 20454 35848 20482
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 35728 20058 35756 20334
rect 35716 20052 35768 20058
rect 35716 19994 35768 20000
rect 35820 19938 35848 20454
rect 35584 18844 35664 18850
rect 35532 18838 35664 18844
rect 35544 18822 35664 18838
rect 35728 19910 35848 19938
rect 35624 18760 35676 18766
rect 35624 18702 35676 18708
rect 35440 18624 35492 18630
rect 35440 18566 35492 18572
rect 35348 17876 35400 17882
rect 35348 17818 35400 17824
rect 35452 17814 35480 18566
rect 35256 17808 35308 17814
rect 35256 17750 35308 17756
rect 35440 17808 35492 17814
rect 35440 17750 35492 17756
rect 35268 17678 35296 17750
rect 35256 17672 35308 17678
rect 35256 17614 35308 17620
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 34888 17536 34940 17542
rect 34888 17478 34940 17484
rect 34900 17338 34928 17478
rect 34888 17332 34940 17338
rect 34888 17274 34940 17280
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34704 16788 34756 16794
rect 34704 16730 34756 16736
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 35360 16658 35388 16730
rect 34704 16652 34756 16658
rect 34704 16594 34756 16600
rect 35348 16652 35400 16658
rect 35348 16594 35400 16600
rect 34520 16584 34572 16590
rect 34520 16526 34572 16532
rect 34532 16182 34560 16526
rect 34520 16176 34572 16182
rect 34520 16118 34572 16124
rect 34336 15904 34388 15910
rect 34336 15846 34388 15852
rect 34348 15570 34376 15846
rect 34336 15564 34388 15570
rect 34336 15506 34388 15512
rect 34532 15366 34560 16118
rect 34716 15978 34744 16594
rect 34796 16448 34848 16454
rect 34796 16390 34848 16396
rect 34808 16250 34836 16390
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 34796 16108 34848 16114
rect 34796 16050 34848 16056
rect 34704 15972 34756 15978
rect 34704 15914 34756 15920
rect 34808 15706 34836 16050
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 35254 15600 35310 15609
rect 35254 15535 35256 15544
rect 35308 15535 35310 15544
rect 35256 15506 35308 15512
rect 34704 15428 34756 15434
rect 34704 15370 34756 15376
rect 34520 15360 34572 15366
rect 34520 15302 34572 15308
rect 34428 15020 34480 15026
rect 34428 14962 34480 14968
rect 34440 12442 34468 14962
rect 34612 14544 34664 14550
rect 34612 14486 34664 14492
rect 34520 13184 34572 13190
rect 34520 13126 34572 13132
rect 34532 12918 34560 13126
rect 34520 12912 34572 12918
rect 34520 12854 34572 12860
rect 34624 12782 34652 14486
rect 34612 12776 34664 12782
rect 34612 12718 34664 12724
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34428 12436 34480 12442
rect 34428 12378 34480 12384
rect 34624 11830 34652 12582
rect 34612 11824 34664 11830
rect 34612 11766 34664 11772
rect 34716 11286 34744 15370
rect 34796 15360 34848 15366
rect 34796 15302 34848 15308
rect 35256 15360 35308 15366
rect 35256 15302 35308 15308
rect 34808 15094 34836 15302
rect 34796 15088 34848 15094
rect 34796 15030 34848 15036
rect 34808 13326 34836 15030
rect 35268 14890 35296 15302
rect 35360 14958 35388 16594
rect 35544 16266 35572 17614
rect 35636 16946 35664 18702
rect 35728 17134 35756 19910
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 35808 19304 35860 19310
rect 35808 19246 35860 19252
rect 35820 17678 35848 19246
rect 35912 18970 35940 19382
rect 35900 18964 35952 18970
rect 35900 18906 35952 18912
rect 35900 18828 35952 18834
rect 35900 18770 35952 18776
rect 35912 18358 35940 18770
rect 36004 18766 36032 20488
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 35900 18352 35952 18358
rect 35900 18294 35952 18300
rect 36188 18290 36216 22918
rect 36556 22574 36584 23462
rect 36544 22568 36596 22574
rect 36728 22568 36780 22574
rect 36544 22510 36596 22516
rect 36726 22536 36728 22545
rect 36780 22536 36782 22545
rect 36452 22500 36504 22506
rect 36726 22471 36782 22480
rect 36452 22442 36504 22448
rect 36464 21010 36492 22442
rect 36452 21004 36504 21010
rect 36452 20946 36504 20952
rect 36728 20800 36780 20806
rect 36728 20742 36780 20748
rect 36544 20528 36596 20534
rect 36544 20470 36596 20476
rect 36556 19514 36584 20470
rect 36740 19514 36768 20742
rect 36544 19508 36596 19514
rect 36544 19450 36596 19456
rect 36728 19508 36780 19514
rect 36728 19450 36780 19456
rect 36556 18902 36584 19450
rect 36544 18896 36596 18902
rect 36544 18838 36596 18844
rect 36360 18692 36412 18698
rect 36360 18634 36412 18640
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 36176 18284 36228 18290
rect 36176 18226 36228 18232
rect 35808 17672 35860 17678
rect 35808 17614 35860 17620
rect 35716 17128 35768 17134
rect 35716 17070 35768 17076
rect 35636 16918 35848 16946
rect 35544 16238 35756 16266
rect 35532 16176 35584 16182
rect 35532 16118 35584 16124
rect 35440 15496 35492 15502
rect 35440 15438 35492 15444
rect 35452 15026 35480 15438
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35348 14952 35400 14958
rect 35348 14894 35400 14900
rect 35256 14884 35308 14890
rect 35256 14826 35308 14832
rect 35348 14816 35400 14822
rect 35348 14758 35400 14764
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 35360 14550 35388 14758
rect 35348 14544 35400 14550
rect 35348 14486 35400 14492
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 35176 13841 35204 14282
rect 35452 14090 35480 14962
rect 35360 14062 35480 14090
rect 35162 13832 35218 13841
rect 35162 13767 35218 13776
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 35360 13512 35388 14062
rect 35440 14000 35492 14006
rect 35440 13942 35492 13948
rect 35268 13484 35388 13512
rect 35164 13456 35216 13462
rect 35164 13398 35216 13404
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 35176 13258 35204 13398
rect 35268 13326 35296 13484
rect 35256 13320 35308 13326
rect 35256 13262 35308 13268
rect 35164 13252 35216 13258
rect 35164 13194 35216 13200
rect 35348 13184 35400 13190
rect 35348 13126 35400 13132
rect 35360 12850 35388 13126
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35348 11824 35400 11830
rect 35348 11766 35400 11772
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34704 11280 34756 11286
rect 34704 11222 34756 11228
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 35360 10266 35388 11766
rect 35452 11354 35480 13942
rect 35544 12434 35572 16118
rect 35728 15910 35756 16238
rect 35716 15904 35768 15910
rect 35716 15846 35768 15852
rect 35624 15496 35676 15502
rect 35624 15438 35676 15444
rect 35636 15094 35664 15438
rect 35728 15366 35756 15846
rect 35716 15360 35768 15366
rect 35716 15302 35768 15308
rect 35624 15088 35676 15094
rect 35624 15030 35676 15036
rect 35820 15026 35848 16918
rect 35900 16652 35952 16658
rect 35900 16594 35952 16600
rect 35716 15020 35768 15026
rect 35716 14962 35768 14968
rect 35808 15020 35860 15026
rect 35808 14962 35860 14968
rect 35728 14074 35756 14962
rect 35808 14816 35860 14822
rect 35808 14758 35860 14764
rect 35716 14068 35768 14074
rect 35636 14028 35716 14056
rect 35636 13394 35664 14028
rect 35716 14010 35768 14016
rect 35716 13864 35768 13870
rect 35716 13806 35768 13812
rect 35624 13388 35676 13394
rect 35624 13330 35676 13336
rect 35728 12918 35756 13806
rect 35716 12912 35768 12918
rect 35716 12854 35768 12860
rect 35820 12850 35848 14758
rect 35808 12844 35860 12850
rect 35808 12786 35860 12792
rect 35624 12436 35676 12442
rect 35544 12406 35624 12434
rect 35624 12378 35676 12384
rect 35912 11558 35940 16594
rect 35992 13320 36044 13326
rect 35992 13262 36044 13268
rect 35900 11552 35952 11558
rect 35900 11494 35952 11500
rect 35440 11348 35492 11354
rect 35440 11290 35492 11296
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35348 10260 35400 10266
rect 35348 10202 35400 10208
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 35452 9178 35480 11154
rect 35624 11076 35676 11082
rect 35624 11018 35676 11024
rect 35636 10266 35664 11018
rect 35806 10976 35862 10985
rect 35806 10911 35862 10920
rect 35820 10606 35848 10911
rect 35808 10600 35860 10606
rect 35808 10542 35860 10548
rect 35624 10260 35676 10266
rect 35624 10202 35676 10208
rect 36004 9586 36032 13262
rect 36096 12918 36124 18226
rect 36268 18080 36320 18086
rect 36268 18022 36320 18028
rect 36280 17202 36308 18022
rect 36268 17196 36320 17202
rect 36268 17138 36320 17144
rect 36280 16522 36308 17138
rect 36268 16516 36320 16522
rect 36268 16458 36320 16464
rect 36372 15094 36400 18634
rect 36556 16046 36584 18838
rect 36740 18426 36768 19450
rect 36728 18420 36780 18426
rect 36728 18362 36780 18368
rect 36636 18080 36688 18086
rect 36636 18022 36688 18028
rect 36544 16040 36596 16046
rect 36544 15982 36596 15988
rect 36556 15162 36584 15982
rect 36544 15156 36596 15162
rect 36544 15098 36596 15104
rect 36360 15088 36412 15094
rect 36360 15030 36412 15036
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 36084 12912 36136 12918
rect 36084 12854 36136 12860
rect 36084 12776 36136 12782
rect 36084 12718 36136 12724
rect 36096 11898 36124 12718
rect 36084 11892 36136 11898
rect 36084 11834 36136 11840
rect 36084 11280 36136 11286
rect 36084 11222 36136 11228
rect 36096 11150 36124 11222
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 36188 9518 36216 14350
rect 36556 14006 36584 15098
rect 36544 14000 36596 14006
rect 36544 13942 36596 13948
rect 36452 13864 36504 13870
rect 36452 13806 36504 13812
rect 36268 13184 36320 13190
rect 36268 13126 36320 13132
rect 36280 12782 36308 13126
rect 36464 12986 36492 13806
rect 36452 12980 36504 12986
rect 36452 12922 36504 12928
rect 36648 12850 36676 18022
rect 36728 17128 36780 17134
rect 36726 17096 36728 17105
rect 36780 17096 36782 17105
rect 36726 17031 36782 17040
rect 36728 14816 36780 14822
rect 36728 14758 36780 14764
rect 36740 14482 36768 14758
rect 36728 14476 36780 14482
rect 36728 14418 36780 14424
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 36268 12776 36320 12782
rect 36268 12718 36320 12724
rect 36648 12434 36676 12786
rect 36648 12406 36860 12434
rect 36832 12306 36860 12406
rect 36820 12300 36872 12306
rect 36820 12242 36872 12248
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 36176 9512 36228 9518
rect 36176 9454 36228 9460
rect 36280 9450 36308 12174
rect 36726 11792 36782 11801
rect 36726 11727 36728 11736
rect 36780 11727 36782 11736
rect 36728 11698 36780 11704
rect 36544 11552 36596 11558
rect 36544 11494 36596 11500
rect 36556 10742 36584 11494
rect 36832 11286 36860 12242
rect 36820 11280 36872 11286
rect 36820 11222 36872 11228
rect 36636 11076 36688 11082
rect 36636 11018 36688 11024
rect 36544 10736 36596 10742
rect 36544 10678 36596 10684
rect 36452 10464 36504 10470
rect 36452 10406 36504 10412
rect 36464 10130 36492 10406
rect 36452 10124 36504 10130
rect 36452 10066 36504 10072
rect 36648 9654 36676 11018
rect 36728 10600 36780 10606
rect 36728 10542 36780 10548
rect 36636 9648 36688 9654
rect 36636 9590 36688 9596
rect 36268 9444 36320 9450
rect 36268 9386 36320 9392
rect 35440 9172 35492 9178
rect 35440 9114 35492 9120
rect 36740 8498 36768 10542
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35636 7410 35664 7822
rect 35624 7404 35676 7410
rect 35624 7346 35676 7352
rect 36268 7200 36320 7206
rect 36268 7142 36320 7148
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34256 6886 34468 6914
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 28816 6316 28868 6322
rect 28816 6258 28868 6264
rect 30392 5710 30420 6734
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 26424 5160 26476 5166
rect 26424 5102 26476 5108
rect 28264 5160 28316 5166
rect 28264 5102 28316 5108
rect 26436 4690 26464 5102
rect 32588 5024 32640 5030
rect 32588 4966 32640 4972
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 25964 4548 26016 4554
rect 25964 4490 26016 4496
rect 26240 4548 26292 4554
rect 26240 4490 26292 4496
rect 25780 4480 25832 4486
rect 25780 4422 25832 4428
rect 25792 4146 25820 4422
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 24674 4040 24730 4049
rect 24674 3975 24730 3984
rect 24688 3534 24716 3975
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31390 3904 31446 3913
rect 31220 3602 31248 3878
rect 31390 3839 31446 3848
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21376 2746 21588 2774
rect 21560 2378 21588 2746
rect 21548 2372 21600 2378
rect 21548 2314 21600 2320
rect 21192 1686 21312 1714
rect 21284 800 21312 1686
rect 21928 800 21956 2790
rect 22020 2650 22048 2926
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 22480 2650 22508 2858
rect 22572 2650 22600 3470
rect 24308 3460 24360 3466
rect 24308 3402 24360 3408
rect 30748 3460 30800 3466
rect 30748 3402 30800 3408
rect 24320 3126 24348 3402
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 3126 24808 3334
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 30760 3058 30788 3402
rect 31404 3058 31432 3839
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 30748 3052 30800 3058
rect 30748 2994 30800 3000
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24596 2650 24624 2926
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 25148 800 25176 2926
rect 31588 800 31616 3538
rect 31772 2582 31800 4558
rect 32404 4548 32456 4554
rect 32404 4490 32456 4496
rect 32416 3194 32444 4490
rect 32600 4146 32628 4966
rect 33140 4684 33192 4690
rect 33140 4626 33192 4632
rect 32588 4140 32640 4146
rect 32588 4082 32640 4088
rect 32496 3664 32548 3670
rect 32496 3606 32548 3612
rect 32508 3194 32536 3606
rect 32404 3188 32456 3194
rect 32404 3130 32456 3136
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 32140 2650 32168 2926
rect 32220 2916 32272 2922
rect 32220 2858 32272 2864
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 31760 2576 31812 2582
rect 31760 2518 31812 2524
rect 32232 800 32260 2858
rect 33152 2802 33180 4626
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 33508 4072 33560 4078
rect 33508 4014 33560 4020
rect 33428 3738 33456 4014
rect 33416 3732 33468 3738
rect 33416 3674 33468 3680
rect 32876 2774 33180 2802
rect 32876 800 32904 2774
rect 33520 800 33548 4014
rect 33600 3936 33652 3942
rect 33600 3878 33652 3884
rect 33612 3534 33640 3878
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34440 3466 34468 6886
rect 36280 6866 36308 7142
rect 36268 6860 36320 6866
rect 36268 6802 36320 6808
rect 36452 6724 36504 6730
rect 36452 6666 36504 6672
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 34440 2854 34468 3402
rect 34428 2848 34480 2854
rect 34428 2790 34480 2796
rect 34532 2446 34560 5646
rect 36464 5370 36492 6666
rect 36728 6112 36780 6118
rect 36728 6054 36780 6060
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36634 5264 36690 5273
rect 36634 5199 36636 5208
rect 36688 5199 36690 5208
rect 36636 5170 36688 5176
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 36636 5024 36688 5030
rect 36636 4966 36688 4972
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 34716 3534 34744 4558
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34808 3058 34836 4966
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35808 4072 35860 4078
rect 35808 4014 35860 4020
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35072 3392 35124 3398
rect 35072 3334 35124 3340
rect 35084 3126 35112 3334
rect 35072 3120 35124 3126
rect 35072 3062 35124 3068
rect 34796 3052 34848 3058
rect 34796 2994 34848 3000
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34520 2440 34572 2446
rect 34520 2382 34572 2388
rect 35164 2372 35216 2378
rect 35164 2314 35216 2320
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35176 105 35204 2314
rect 35452 800 35480 2926
rect 35820 2145 35848 4014
rect 36648 3754 36676 4966
rect 36740 4146 36768 6054
rect 36728 4140 36780 4146
rect 36728 4082 36780 4088
rect 36648 3726 36768 3754
rect 36544 2848 36596 2854
rect 36544 2790 36596 2796
rect 36556 2514 36584 2790
rect 36740 2514 36768 3726
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 36544 2508 36596 2514
rect 36544 2450 36596 2456
rect 36728 2508 36780 2514
rect 36728 2450 36780 2456
rect 35806 2136 35862 2145
rect 35806 2071 35862 2080
rect 36832 1714 36860 3538
rect 36924 2446 36952 30874
rect 37186 29336 37242 29345
rect 37186 29271 37242 29280
rect 37200 28626 37228 29271
rect 37188 28620 37240 28626
rect 37188 28562 37240 28568
rect 37292 26330 37320 37198
rect 37384 34066 37412 39200
rect 37924 37256 37976 37262
rect 37924 37198 37976 37204
rect 37464 36100 37516 36106
rect 37464 36042 37516 36048
rect 37476 35834 37504 36042
rect 37464 35828 37516 35834
rect 37464 35770 37516 35776
rect 37936 35290 37964 37198
rect 38028 35766 38056 39200
rect 38106 36816 38162 36825
rect 38106 36751 38162 36760
rect 38568 36780 38620 36786
rect 38120 36242 38148 36751
rect 38568 36722 38620 36728
rect 38108 36236 38160 36242
rect 38108 36178 38160 36184
rect 38016 35760 38068 35766
rect 38016 35702 38068 35708
rect 38384 35692 38436 35698
rect 38384 35634 38436 35640
rect 38016 35488 38068 35494
rect 38016 35430 38068 35436
rect 37924 35284 37976 35290
rect 37924 35226 37976 35232
rect 37556 35012 37608 35018
rect 37556 34954 37608 34960
rect 37568 34746 37596 34954
rect 37556 34740 37608 34746
rect 37556 34682 37608 34688
rect 37372 34060 37424 34066
rect 37372 34002 37424 34008
rect 37372 33924 37424 33930
rect 37372 33866 37424 33872
rect 37384 33658 37412 33866
rect 37372 33652 37424 33658
rect 37372 33594 37424 33600
rect 37556 33448 37608 33454
rect 37556 33390 37608 33396
rect 37568 30258 37596 33390
rect 37648 32836 37700 32842
rect 37648 32778 37700 32784
rect 37660 32570 37688 32778
rect 37648 32564 37700 32570
rect 37648 32506 37700 32512
rect 37936 32434 37964 35226
rect 37924 32428 37976 32434
rect 37924 32370 37976 32376
rect 37936 31346 37964 32370
rect 37924 31340 37976 31346
rect 37924 31282 37976 31288
rect 37556 30252 37608 30258
rect 37608 30212 37780 30240
rect 37556 30194 37608 30200
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37476 29714 37504 29990
rect 37464 29708 37516 29714
rect 37464 29650 37516 29656
rect 37554 29200 37610 29209
rect 37554 29135 37556 29144
rect 37608 29135 37610 29144
rect 37556 29106 37608 29112
rect 37372 27396 37424 27402
rect 37372 27338 37424 27344
rect 37384 27130 37412 27338
rect 37372 27124 37424 27130
rect 37372 27066 37424 27072
rect 37464 26988 37516 26994
rect 37464 26930 37516 26936
rect 37292 26302 37412 26330
rect 37280 26240 37332 26246
rect 37280 26182 37332 26188
rect 37292 25906 37320 26182
rect 37280 25900 37332 25906
rect 37280 25842 37332 25848
rect 37384 25786 37412 26302
rect 37292 25758 37412 25786
rect 37292 24682 37320 25758
rect 37280 24676 37332 24682
rect 37280 24618 37332 24624
rect 37292 23730 37320 24618
rect 37372 24132 37424 24138
rect 37372 24074 37424 24080
rect 37384 23866 37412 24074
rect 37372 23860 37424 23866
rect 37372 23802 37424 23808
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37476 23662 37504 26930
rect 37464 23656 37516 23662
rect 37464 23598 37516 23604
rect 37476 22642 37504 23598
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37004 22568 37056 22574
rect 37004 22510 37056 22516
rect 37016 9586 37044 22510
rect 37280 22432 37332 22438
rect 37280 22374 37332 22380
rect 37188 22228 37240 22234
rect 37188 22170 37240 22176
rect 37094 20496 37150 20505
rect 37094 20431 37150 20440
rect 37108 19922 37136 20431
rect 37096 19916 37148 19922
rect 37096 19858 37148 19864
rect 37094 18456 37150 18465
rect 37094 18391 37150 18400
rect 37108 17746 37136 18391
rect 37096 17740 37148 17746
rect 37096 17682 37148 17688
rect 37096 15564 37148 15570
rect 37096 15506 37148 15512
rect 37108 14385 37136 15506
rect 37094 14376 37150 14385
rect 37094 14311 37150 14320
rect 37200 12434 37228 22170
rect 37292 22094 37320 22374
rect 37292 22066 37412 22094
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37292 21350 37320 21898
rect 37280 21344 37332 21350
rect 37280 21286 37332 21292
rect 37292 20874 37320 21286
rect 37280 20868 37332 20874
rect 37280 20810 37332 20816
rect 37292 20534 37320 20810
rect 37280 20528 37332 20534
rect 37280 20470 37332 20476
rect 37384 20330 37412 22066
rect 37464 22092 37516 22098
rect 37464 22034 37516 22040
rect 37476 21865 37504 22034
rect 37462 21856 37518 21865
rect 37462 21791 37518 21800
rect 37568 21554 37596 29106
rect 37648 25900 37700 25906
rect 37648 25842 37700 25848
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37372 20324 37424 20330
rect 37372 20266 37424 20272
rect 37372 19712 37424 19718
rect 37372 19654 37424 19660
rect 37384 19446 37412 19654
rect 37372 19440 37424 19446
rect 37372 19382 37424 19388
rect 37476 19378 37504 20402
rect 37464 19372 37516 19378
rect 37464 19314 37516 19320
rect 37476 17814 37504 19314
rect 37464 17808 37516 17814
rect 37464 17750 37516 17756
rect 37464 16720 37516 16726
rect 37464 16662 37516 16668
rect 37476 16114 37504 16662
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37464 14612 37516 14618
rect 37464 14554 37516 14560
rect 37476 13938 37504 14554
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 37108 12406 37228 12434
rect 37004 9580 37056 9586
rect 37004 9522 37056 9528
rect 37108 6390 37136 12406
rect 37186 9616 37242 9625
rect 37186 9551 37242 9560
rect 37200 9042 37228 9551
rect 37188 9036 37240 9042
rect 37188 8978 37240 8984
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 37096 6384 37148 6390
rect 37096 6326 37148 6332
rect 37096 5772 37148 5778
rect 37096 5714 37148 5720
rect 36912 2440 36964 2446
rect 36912 2382 36964 2388
rect 36740 1686 36860 1714
rect 36740 800 36768 1686
rect 35162 96 35218 105
rect 35162 31 35218 40
rect 35410 0 35522 800
rect 36698 0 36810 800
rect 37108 785 37136 5714
rect 37200 5545 37228 6802
rect 37186 5536 37242 5545
rect 37186 5471 37242 5480
rect 37280 4684 37332 4690
rect 37280 4626 37332 4632
rect 37292 4146 37320 4626
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 37372 3460 37424 3466
rect 37372 3402 37424 3408
rect 37384 800 37412 3402
rect 37476 3058 37504 13874
rect 37568 12850 37596 21490
rect 37660 18850 37688 25842
rect 37752 19122 37780 30212
rect 37924 28960 37976 28966
rect 37924 28902 37976 28908
rect 37936 28626 37964 28902
rect 37924 28620 37976 28626
rect 37924 28562 37976 28568
rect 37924 26376 37976 26382
rect 37924 26318 37976 26324
rect 37832 24608 37884 24614
rect 37832 24550 37884 24556
rect 37844 19990 37872 24550
rect 37936 23066 37964 26318
rect 38028 23186 38056 35430
rect 38108 35080 38160 35086
rect 38108 35022 38160 35028
rect 38120 33522 38148 35022
rect 38292 34604 38344 34610
rect 38292 34546 38344 34552
rect 38108 33516 38160 33522
rect 38108 33458 38160 33464
rect 38108 32836 38160 32842
rect 38108 32778 38160 32784
rect 38120 32745 38148 32778
rect 38106 32736 38162 32745
rect 38106 32671 38162 32680
rect 38108 31816 38160 31822
rect 38108 31758 38160 31764
rect 38120 31385 38148 31758
rect 38106 31376 38162 31385
rect 38106 31311 38162 31320
rect 38106 30696 38162 30705
rect 38106 30631 38108 30640
rect 38160 30631 38162 30640
rect 38108 30602 38160 30608
rect 38106 30016 38162 30025
rect 38106 29951 38162 29960
rect 38120 29714 38148 29951
rect 38108 29708 38160 29714
rect 38108 29650 38160 29656
rect 38108 28552 38160 28558
rect 38108 28494 38160 28500
rect 38120 28082 38148 28494
rect 38108 28076 38160 28082
rect 38108 28018 38160 28024
rect 38106 25936 38162 25945
rect 38106 25871 38162 25880
rect 38120 25362 38148 25871
rect 38200 25696 38252 25702
rect 38200 25638 38252 25644
rect 38108 25356 38160 25362
rect 38108 25298 38160 25304
rect 38108 24132 38160 24138
rect 38108 24074 38160 24080
rect 38120 23905 38148 24074
rect 38106 23896 38162 23905
rect 38106 23831 38162 23840
rect 38016 23180 38068 23186
rect 38016 23122 38068 23128
rect 37936 23038 38056 23066
rect 37924 22432 37976 22438
rect 37924 22374 37976 22380
rect 37936 22098 37964 22374
rect 37924 22092 37976 22098
rect 37924 22034 37976 22040
rect 37924 21344 37976 21350
rect 37924 21286 37976 21292
rect 37832 19984 37884 19990
rect 37832 19926 37884 19932
rect 37936 19922 37964 21286
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 37752 19094 37872 19122
rect 37660 18822 37780 18850
rect 37648 18692 37700 18698
rect 37648 18634 37700 18640
rect 37660 18426 37688 18634
rect 37648 18420 37700 18426
rect 37648 18362 37700 18368
rect 37648 13252 37700 13258
rect 37648 13194 37700 13200
rect 37660 12986 37688 13194
rect 37648 12980 37700 12986
rect 37648 12922 37700 12928
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37752 12434 37780 18822
rect 37844 16114 37872 19094
rect 37924 18080 37976 18086
rect 37924 18022 37976 18028
rect 37936 17746 37964 18022
rect 38028 17814 38056 23038
rect 38212 22098 38240 25638
rect 38200 22092 38252 22098
rect 38200 22034 38252 22040
rect 38106 21176 38162 21185
rect 38106 21111 38162 21120
rect 38120 21010 38148 21111
rect 38108 21004 38160 21010
rect 38108 20946 38160 20952
rect 38016 17808 38068 17814
rect 38016 17750 38068 17756
rect 37924 17740 37976 17746
rect 37924 17682 37976 17688
rect 37924 16516 37976 16522
rect 37924 16458 37976 16464
rect 38108 16516 38160 16522
rect 38108 16458 38160 16464
rect 37936 16250 37964 16458
rect 38120 16425 38148 16458
rect 38106 16416 38162 16425
rect 38106 16351 38162 16360
rect 37924 16244 37976 16250
rect 37924 16186 37976 16192
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 38108 15496 38160 15502
rect 38108 15438 38160 15444
rect 37924 15428 37976 15434
rect 37924 15370 37976 15376
rect 37936 14074 37964 15370
rect 38120 15178 38148 15438
rect 38028 15150 38148 15178
rect 37924 14068 37976 14074
rect 37924 14010 37976 14016
rect 37752 12406 37872 12434
rect 37648 12164 37700 12170
rect 37648 12106 37700 12112
rect 37660 11898 37688 12106
rect 37648 11892 37700 11898
rect 37648 11834 37700 11840
rect 37740 11756 37792 11762
rect 37740 11698 37792 11704
rect 37556 4548 37608 4554
rect 37556 4490 37608 4496
rect 37568 4185 37596 4490
rect 37554 4176 37610 4185
rect 37554 4111 37610 4120
rect 37752 3534 37780 11698
rect 37844 4162 37872 12406
rect 37924 9376 37976 9382
rect 37924 9318 37976 9324
rect 37936 9042 37964 9318
rect 37924 9036 37976 9042
rect 37924 8978 37976 8984
rect 38028 8090 38056 15150
rect 38106 15056 38162 15065
rect 38304 15026 38332 34546
rect 38106 14991 38162 15000
rect 38292 15020 38344 15026
rect 38120 14482 38148 14991
rect 38292 14962 38344 14968
rect 38108 14476 38160 14482
rect 38108 14418 38160 14424
rect 38106 13696 38162 13705
rect 38106 13631 38162 13640
rect 38120 13394 38148 13631
rect 38108 13388 38160 13394
rect 38108 13330 38160 13336
rect 38108 12164 38160 12170
rect 38108 12106 38160 12112
rect 38120 11665 38148 12106
rect 38106 11656 38162 11665
rect 38106 11591 38162 11600
rect 38200 11076 38252 11082
rect 38200 11018 38252 11024
rect 38106 10296 38162 10305
rect 38106 10231 38162 10240
rect 38120 10130 38148 10231
rect 38108 10124 38160 10130
rect 38108 10066 38160 10072
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 38120 8498 38148 8910
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38016 8084 38068 8090
rect 38016 8026 38068 8032
rect 38016 6316 38068 6322
rect 38016 6258 38068 6264
rect 38028 6225 38056 6258
rect 38014 6216 38070 6225
rect 38014 6151 38070 6160
rect 38108 5704 38160 5710
rect 38108 5646 38160 5652
rect 37924 5636 37976 5642
rect 37924 5578 37976 5584
rect 37936 5370 37964 5578
rect 37924 5364 37976 5370
rect 37924 5306 37976 5312
rect 37844 4134 37964 4162
rect 38120 4146 38148 5646
rect 37832 4072 37884 4078
rect 37832 4014 37884 4020
rect 37844 3738 37872 4014
rect 37936 3942 37964 4134
rect 38108 4140 38160 4146
rect 38108 4082 38160 4088
rect 37924 3936 37976 3942
rect 37924 3878 37976 3884
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 37924 3664 37976 3670
rect 37924 3606 37976 3612
rect 37740 3528 37792 3534
rect 37740 3470 37792 3476
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37936 2650 37964 3606
rect 38212 3466 38240 11018
rect 38396 9586 38424 35634
rect 38580 10674 38608 36722
rect 38658 32056 38714 32065
rect 38658 31991 38714 32000
rect 38672 27538 38700 31991
rect 38660 27532 38712 27538
rect 38660 27474 38712 27480
rect 38568 10668 38620 10674
rect 38568 10610 38620 10616
rect 38384 9580 38436 9586
rect 38384 9522 38436 9528
rect 38660 7812 38712 7818
rect 38660 7754 38712 7760
rect 38200 3460 38252 3466
rect 38200 3402 38252 3408
rect 37924 2644 37976 2650
rect 37924 2586 37976 2592
rect 38016 2576 38068 2582
rect 38016 2518 38068 2524
rect 38028 800 38056 2518
rect 38672 800 38700 7754
rect 37094 776 37150 785
rect 37094 711 37150 720
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
<< via2 >>
rect 1582 37440 1638 37496
rect 2870 38800 2926 38856
rect 1398 36760 1454 36816
rect 1398 32000 1454 32056
rect 2778 36080 2834 36136
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2318 34604 2374 34640
rect 2318 34584 2320 34604
rect 2320 34584 2372 34604
rect 2372 34584 2374 34604
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 3974 34720 4030 34776
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 3422 33380 3478 33416
rect 3422 33360 3424 33380
rect 3424 33360 3476 33380
rect 3476 33360 3478 33380
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 2870 25880 2926 25936
rect 2318 25200 2374 25256
rect 1858 19760 1914 19816
rect 2134 19080 2190 19136
rect 1398 15680 1454 15736
rect 1398 14356 1400 14376
rect 1400 14356 1452 14376
rect 1452 14356 1454 14376
rect 1398 14320 1454 14356
rect 2042 11636 2044 11656
rect 2044 11636 2096 11656
rect 2096 11636 2098 11656
rect 2042 11600 2098 11636
rect 1858 8880 1914 8936
rect 4158 29008 4214 29064
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2778 13640 2834 13696
rect 2778 12300 2834 12336
rect 2778 12280 2780 12300
rect 2780 12280 2832 12300
rect 2832 12280 2834 12300
rect 2778 7520 2834 7576
rect 2778 6196 2780 6216
rect 2780 6196 2832 6216
rect 2832 6196 2834 6216
rect 2778 6160 2834 6196
rect 1766 4800 1822 4856
rect 1398 2080 1454 2136
rect 2778 2760 2834 2816
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3974 8200 4030 8256
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3422 4156 3424 4176
rect 3424 4156 3476 4176
rect 3476 4156 3478 4176
rect 3422 4120 3478 4156
rect 3422 3440 3478 3496
rect 2870 1400 2926 1456
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7194 36780 7250 36816
rect 7194 36760 7196 36780
rect 7196 36760 7248 36780
rect 7248 36760 7250 36780
rect 5722 35672 5778 35728
rect 7470 33924 7526 33960
rect 7470 33904 7472 33924
rect 7472 33904 7524 33924
rect 7524 33904 7526 33924
rect 7194 32952 7250 33008
rect 5446 29008 5502 29064
rect 5170 3984 5226 4040
rect 7194 22072 7250 22128
rect 7838 22072 7894 22128
rect 10230 22072 10286 22128
rect 12622 33768 12678 33824
rect 11886 30540 11888 30560
rect 11888 30540 11940 30560
rect 11940 30540 11942 30560
rect 11886 30504 11942 30540
rect 12254 29416 12310 29472
rect 13634 29416 13690 29472
rect 16302 35536 16358 35592
rect 15566 33768 15622 33824
rect 18510 36760 18566 36816
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 11334 22108 11336 22128
rect 11336 22108 11388 22128
rect 11388 22108 11390 22128
rect 11334 22072 11390 22108
rect 11886 19488 11942 19544
rect 13634 20440 13690 20496
rect 13910 19352 13966 19408
rect 14370 23432 14426 23488
rect 14370 19352 14426 19408
rect 15290 22072 15346 22128
rect 15106 19760 15162 19816
rect 15014 19488 15070 19544
rect 16762 30504 16818 30560
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19522 35692 19578 35728
rect 19522 35672 19524 35692
rect 19524 35672 19576 35692
rect 19576 35672 19578 35692
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 20810 35572 20812 35592
rect 20812 35572 20864 35592
rect 20864 35572 20866 35592
rect 20810 35536 20866 35572
rect 21454 32952 21510 33008
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 16762 19508 16818 19544
rect 16762 19488 16764 19508
rect 16764 19488 16816 19508
rect 16816 19488 16818 19508
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 17866 20440 17922 20496
rect 17314 19760 17370 19816
rect 18418 19352 18474 19408
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 18602 19488 18658 19544
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20534 22480 20590 22536
rect 21270 25200 21326 25256
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19246 16632 19302 16688
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20718 20032 20774 20088
rect 20718 19760 20774 19816
rect 19062 12416 19118 12472
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19338 9968 19394 10024
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20074 8880 20130 8936
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19430 7248 19486 7304
rect 21178 23160 21234 23216
rect 20258 8880 20314 8936
rect 20902 14612 20958 14648
rect 20902 14592 20904 14612
rect 20904 14592 20956 14612
rect 20956 14592 20958 14612
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 21454 22208 21510 22264
rect 22374 35944 22430 36000
rect 24582 33904 24638 33960
rect 23570 26852 23626 26888
rect 23570 26832 23572 26852
rect 23572 26832 23624 26852
rect 23624 26832 23626 26852
rect 21086 7792 21142 7848
rect 20902 7520 20958 7576
rect 20718 3984 20774 4040
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22374 19896 22430 19952
rect 21546 10784 21602 10840
rect 21454 7964 21456 7984
rect 21456 7964 21508 7984
rect 21508 7964 21510 7984
rect 21454 7928 21510 7964
rect 23018 22380 23020 22400
rect 23020 22380 23072 22400
rect 23072 22380 23074 22400
rect 23018 22344 23074 22380
rect 23018 19252 23020 19272
rect 23020 19252 23072 19272
rect 23072 19252 23074 19272
rect 23018 19216 23074 19252
rect 25502 29280 25558 29336
rect 23938 21936 23994 21992
rect 23202 16532 23204 16552
rect 23204 16532 23256 16552
rect 23256 16532 23258 16552
rect 23202 16496 23258 16532
rect 22282 8916 22284 8936
rect 22284 8916 22336 8936
rect 22336 8916 22338 8936
rect 22282 8880 22338 8916
rect 26054 29008 26110 29064
rect 26974 29844 27030 29880
rect 26974 29824 26976 29844
rect 26976 29824 27028 29844
rect 27028 29824 27030 29844
rect 27250 30268 27252 30288
rect 27252 30268 27304 30288
rect 27304 30268 27306 30288
rect 27250 30232 27306 30268
rect 27710 30268 27712 30288
rect 27712 30268 27764 30288
rect 27764 30268 27766 30288
rect 27710 30232 27766 30268
rect 37186 38800 37242 38856
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 36726 37440 36782 37496
rect 28078 29824 28134 29880
rect 26330 27412 26332 27432
rect 26332 27412 26384 27432
rect 26384 27412 26386 27432
rect 26330 27376 26386 27412
rect 27342 27548 27344 27568
rect 27344 27548 27396 27568
rect 27396 27548 27398 27568
rect 27342 27512 27398 27548
rect 27434 27240 27490 27296
rect 27894 27376 27950 27432
rect 28446 29300 28502 29336
rect 28446 29280 28448 29300
rect 28448 29280 28500 29300
rect 28500 29280 28502 29300
rect 28170 27532 28226 27568
rect 28170 27512 28172 27532
rect 28172 27512 28224 27532
rect 28224 27512 28226 27532
rect 28354 27240 28410 27296
rect 29734 32444 29736 32464
rect 29736 32444 29788 32464
rect 29788 32444 29790 32464
rect 29734 32408 29790 32444
rect 30470 32816 30526 32872
rect 30746 32000 30802 32056
rect 30746 30368 30802 30424
rect 31298 32852 31300 32872
rect 31300 32852 31352 32872
rect 31352 32852 31354 32872
rect 31298 32816 31354 32852
rect 31666 32444 31668 32464
rect 31668 32444 31720 32464
rect 31720 32444 31722 32464
rect 31666 32408 31722 32444
rect 31942 32816 31998 32872
rect 31482 32000 31538 32056
rect 30378 29008 30434 29064
rect 28446 23160 28502 23216
rect 25134 20324 25190 20360
rect 25134 20304 25136 20324
rect 25136 20304 25188 20324
rect 25188 20304 25190 20324
rect 26146 20304 26202 20360
rect 24214 16108 24270 16144
rect 24214 16088 24216 16108
rect 24216 16088 24268 16108
rect 24268 16088 24270 16108
rect 23662 12280 23718 12336
rect 23662 11056 23718 11112
rect 23662 7248 23718 7304
rect 24122 10784 24178 10840
rect 27434 20460 27490 20496
rect 27434 20440 27436 20460
rect 27436 20440 27488 20460
rect 27488 20440 27490 20460
rect 27894 20304 27950 20360
rect 27618 19216 27674 19272
rect 27250 17992 27306 18048
rect 28262 20476 28264 20496
rect 28264 20476 28316 20496
rect 28316 20476 28318 20496
rect 28262 20440 28318 20476
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 28262 20304 28318 20360
rect 28906 20304 28962 20360
rect 28906 19916 28962 19952
rect 28906 19896 28908 19916
rect 28908 19896 28960 19916
rect 28960 19896 28962 19916
rect 27250 16632 27306 16688
rect 27066 16088 27122 16144
rect 24766 8900 24822 8936
rect 24766 8880 24768 8900
rect 24768 8880 24820 8900
rect 24820 8880 24822 8900
rect 24214 7248 24270 7304
rect 25594 8744 25650 8800
rect 26146 8880 26202 8936
rect 26514 9968 26570 10024
rect 27342 12280 27398 12336
rect 28630 16652 28686 16688
rect 28630 16632 28632 16652
rect 28632 16632 28684 16652
rect 28684 16632 28686 16652
rect 30010 18808 30066 18864
rect 33782 34584 33838 34640
rect 35806 36080 35862 36136
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 32770 32852 32772 32872
rect 32772 32852 32824 32872
rect 32824 32852 32826 32872
rect 32770 32816 32826 32852
rect 37186 34720 37242 34776
rect 33414 32952 33470 33008
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 31298 20324 31354 20360
rect 31298 20304 31300 20324
rect 31300 20304 31352 20324
rect 31352 20304 31354 20324
rect 26330 6976 26386 7032
rect 27158 7828 27160 7848
rect 27160 7828 27212 7848
rect 27212 7828 27214 7848
rect 27158 7792 27214 7828
rect 27434 7384 27490 7440
rect 30286 12824 30342 12880
rect 31482 19760 31538 19816
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 32034 18808 32090 18864
rect 31942 16496 31998 16552
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 36266 26832 36322 26888
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 33230 17992 33286 18048
rect 30470 12180 30472 12200
rect 30472 12180 30524 12200
rect 30524 12180 30526 12200
rect 30470 12144 30526 12180
rect 27986 8744 28042 8800
rect 27802 7964 27804 7984
rect 27804 7964 27856 7984
rect 27856 7964 27858 7984
rect 27802 7928 27858 7964
rect 32402 12860 32404 12880
rect 32404 12860 32456 12880
rect 32456 12860 32458 12880
rect 32402 12824 32458 12860
rect 32494 12280 32550 12336
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34518 18672 34574 18728
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35990 22480 36046 22536
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34978 19216 35034 19272
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34886 18672 34942 18728
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35438 19116 35440 19136
rect 35440 19116 35492 19136
rect 35492 19116 35494 19136
rect 35438 19080 35494 19116
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35254 15564 35310 15600
rect 35254 15544 35256 15564
rect 35256 15544 35308 15564
rect 35308 15544 35310 15564
rect 36726 22516 36728 22536
rect 36728 22516 36780 22536
rect 36780 22516 36782 22536
rect 36726 22480 36782 22516
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35162 13776 35218 13832
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35806 10920 35862 10976
rect 36726 17076 36728 17096
rect 36728 17076 36780 17096
rect 36780 17076 36782 17096
rect 36726 17040 36782 17076
rect 36726 11756 36782 11792
rect 36726 11736 36728 11756
rect 36728 11736 36780 11756
rect 36780 11736 36782 11756
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 24674 3984 24730 4040
rect 31390 3848 31446 3904
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 36634 5228 36690 5264
rect 36634 5208 36636 5228
rect 36636 5208 36688 5228
rect 36688 5208 36690 5228
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35806 2080 35862 2136
rect 37186 29280 37242 29336
rect 38106 36760 38162 36816
rect 37554 29164 37610 29200
rect 37554 29144 37556 29164
rect 37556 29144 37608 29164
rect 37608 29144 37610 29164
rect 37094 20440 37150 20496
rect 37094 18400 37150 18456
rect 37094 14320 37150 14376
rect 37462 21800 37518 21856
rect 37186 9560 37242 9616
rect 35162 40 35218 96
rect 37186 5480 37242 5536
rect 38106 32680 38162 32736
rect 38106 31320 38162 31376
rect 38106 30660 38162 30696
rect 38106 30640 38108 30660
rect 38108 30640 38160 30660
rect 38160 30640 38162 30660
rect 38106 29960 38162 30016
rect 38106 25880 38162 25936
rect 38106 23840 38162 23896
rect 38106 21120 38162 21176
rect 38106 16360 38162 16416
rect 37554 4120 37610 4176
rect 38106 15000 38162 15056
rect 38106 13640 38162 13696
rect 38106 11600 38162 11656
rect 38106 10240 38162 10296
rect 38014 6160 38070 6216
rect 38658 32000 38714 32056
rect 37094 720 37150 776
<< metal3 >>
rect 0 39388 800 39628
rect 0 38858 800 38948
rect 2865 38858 2931 38861
rect 0 38856 2931 38858
rect 0 38800 2870 38856
rect 2926 38800 2931 38856
rect 0 38798 2931 38800
rect 0 38708 800 38798
rect 2865 38795 2931 38798
rect 37181 38858 37247 38861
rect 39200 38858 40000 38948
rect 37181 38856 40000 38858
rect 37181 38800 37186 38856
rect 37242 38800 40000 38856
rect 37181 38798 40000 38800
rect 37181 38795 37247 38798
rect 39200 38708 40000 38798
rect 39200 38028 40000 38268
rect 0 37498 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 1577 37498 1643 37501
rect 0 37496 1643 37498
rect 0 37440 1582 37496
rect 1638 37440 1643 37496
rect 0 37438 1643 37440
rect 0 37348 800 37438
rect 1577 37435 1643 37438
rect 36721 37498 36787 37501
rect 39200 37498 40000 37588
rect 36721 37496 40000 37498
rect 36721 37440 36726 37496
rect 36782 37440 40000 37496
rect 36721 37438 40000 37440
rect 36721 37435 36787 37438
rect 39200 37348 40000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 1393 36818 1459 36821
rect 7189 36820 7255 36821
rect 7189 36818 7236 36820
rect 0 36816 1459 36818
rect 0 36760 1398 36816
rect 1454 36760 1459 36816
rect 0 36758 1459 36760
rect 7108 36816 7236 36818
rect 7300 36818 7306 36820
rect 18505 36818 18571 36821
rect 7300 36816 18571 36818
rect 7108 36760 7194 36816
rect 7300 36760 18510 36816
rect 18566 36760 18571 36816
rect 7108 36758 7236 36760
rect 0 36668 800 36758
rect 1393 36755 1459 36758
rect 7189 36756 7236 36758
rect 7300 36758 18571 36760
rect 7300 36756 7306 36758
rect 7189 36755 7255 36756
rect 18505 36755 18571 36758
rect 38101 36818 38167 36821
rect 39200 36818 40000 36908
rect 38101 36816 40000 36818
rect 38101 36760 38106 36816
rect 38162 36760 40000 36816
rect 38101 36758 40000 36760
rect 38101 36755 38167 36758
rect 39200 36668 40000 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36228
rect 2773 36138 2839 36141
rect 0 36136 2839 36138
rect 0 36080 2778 36136
rect 2834 36080 2839 36136
rect 0 36078 2839 36080
rect 0 35988 800 36078
rect 2773 36075 2839 36078
rect 35801 36138 35867 36141
rect 39200 36138 40000 36228
rect 35801 36136 40000 36138
rect 35801 36080 35806 36136
rect 35862 36080 40000 36136
rect 35801 36078 40000 36080
rect 35801 36075 35867 36078
rect 22369 36002 22435 36005
rect 30966 36002 30972 36004
rect 22369 36000 30972 36002
rect 22369 35944 22374 36000
rect 22430 35944 30972 36000
rect 22369 35942 30972 35944
rect 22369 35939 22435 35942
rect 30966 35940 30972 35942
rect 31036 35940 31042 36004
rect 39200 35988 40000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 5717 35730 5783 35733
rect 19517 35730 19583 35733
rect 5717 35728 19583 35730
rect 5717 35672 5722 35728
rect 5778 35672 19522 35728
rect 19578 35672 19583 35728
rect 5717 35670 19583 35672
rect 5717 35667 5783 35670
rect 19517 35667 19583 35670
rect 16297 35594 16363 35597
rect 20805 35594 20871 35597
rect 21214 35594 21220 35596
rect 16297 35592 21220 35594
rect 0 35308 800 35548
rect 16297 35536 16302 35592
rect 16358 35536 20810 35592
rect 20866 35536 21220 35592
rect 16297 35534 21220 35536
rect 16297 35531 16363 35534
rect 20805 35531 20871 35534
rect 21214 35532 21220 35534
rect 21284 35532 21290 35596
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 39200 35308 40000 35548
rect 0 34778 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 3969 34778 4035 34781
rect 0 34776 4035 34778
rect 0 34720 3974 34776
rect 4030 34720 4035 34776
rect 0 34718 4035 34720
rect 0 34628 800 34718
rect 3969 34715 4035 34718
rect 37181 34778 37247 34781
rect 39200 34778 40000 34868
rect 37181 34776 40000 34778
rect 37181 34720 37186 34776
rect 37242 34720 40000 34776
rect 37181 34718 40000 34720
rect 37181 34715 37247 34718
rect 2313 34642 2379 34645
rect 33777 34642 33843 34645
rect 2313 34640 33843 34642
rect 2313 34584 2318 34640
rect 2374 34584 33782 34640
rect 33838 34584 33843 34640
rect 39200 34628 40000 34718
rect 2313 34582 33843 34584
rect 2313 34579 2379 34582
rect 33777 34579 33843 34582
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 7465 33962 7531 33965
rect 24577 33962 24643 33965
rect 7465 33960 24643 33962
rect 7465 33904 7470 33960
rect 7526 33904 24582 33960
rect 24638 33904 24643 33960
rect 7465 33902 24643 33904
rect 7465 33899 7531 33902
rect 24577 33899 24643 33902
rect 12617 33826 12683 33829
rect 15561 33826 15627 33829
rect 12617 33824 15627 33826
rect 12617 33768 12622 33824
rect 12678 33768 15566 33824
rect 15622 33768 15627 33824
rect 12617 33766 15627 33768
rect 12617 33763 12683 33766
rect 15561 33763 15627 33766
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 3417 33418 3483 33421
rect 0 33416 3483 33418
rect 0 33360 3422 33416
rect 3478 33360 3483 33416
rect 0 33358 3483 33360
rect 0 33268 800 33358
rect 3417 33355 3483 33358
rect 39200 33268 40000 33508
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 7189 33010 7255 33013
rect 20846 33010 20852 33012
rect 7189 33008 20852 33010
rect 7189 32952 7194 33008
rect 7250 32952 20852 33008
rect 7189 32950 20852 32952
rect 7189 32947 7255 32950
rect 20846 32948 20852 32950
rect 20916 33010 20922 33012
rect 21449 33010 21515 33013
rect 33409 33010 33475 33013
rect 20916 33008 33475 33010
rect 20916 32952 21454 33008
rect 21510 32952 33414 33008
rect 33470 32952 33475 33008
rect 20916 32950 33475 32952
rect 20916 32948 20922 32950
rect 21449 32947 21515 32950
rect 33409 32947 33475 32950
rect 30465 32874 30531 32877
rect 31293 32874 31359 32877
rect 30465 32872 31359 32874
rect 30465 32816 30470 32872
rect 30526 32816 31298 32872
rect 31354 32816 31359 32872
rect 30465 32814 31359 32816
rect 30465 32811 30531 32814
rect 31293 32811 31359 32814
rect 31937 32874 32003 32877
rect 32765 32874 32831 32877
rect 31937 32872 32831 32874
rect 31937 32816 31942 32872
rect 31998 32816 32770 32872
rect 32826 32816 32831 32872
rect 31937 32814 32831 32816
rect 31937 32811 32003 32814
rect 32765 32811 32831 32814
rect 38101 32738 38167 32741
rect 39200 32738 40000 32828
rect 38101 32736 40000 32738
rect 38101 32680 38106 32736
rect 38162 32680 40000 32736
rect 38101 32678 40000 32680
rect 38101 32675 38167 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 39200 32588 40000 32678
rect 29729 32466 29795 32469
rect 31661 32466 31727 32469
rect 29729 32464 31727 32466
rect 29729 32408 29734 32464
rect 29790 32408 31666 32464
rect 31722 32408 31727 32464
rect 29729 32406 31727 32408
rect 29729 32403 29795 32406
rect 31661 32403 31727 32406
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1393 32058 1459 32061
rect 0 32056 1459 32058
rect 0 32000 1398 32056
rect 1454 32000 1459 32056
rect 0 31998 1459 32000
rect 0 31908 800 31998
rect 1393 31995 1459 31998
rect 30741 32058 30807 32061
rect 31477 32058 31543 32061
rect 30741 32056 31543 32058
rect 30741 32000 30746 32056
rect 30802 32000 31482 32056
rect 31538 32000 31543 32056
rect 30741 31998 31543 32000
rect 30741 31995 30807 31998
rect 31477 31995 31543 31998
rect 38653 32058 38719 32061
rect 39200 32058 40000 32148
rect 38653 32056 40000 32058
rect 38653 32000 38658 32056
rect 38714 32000 40000 32056
rect 38653 31998 40000 32000
rect 38653 31995 38719 31998
rect 39200 31908 40000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31228 800 31468
rect 38101 31378 38167 31381
rect 39200 31378 40000 31468
rect 38101 31376 40000 31378
rect 38101 31320 38106 31376
rect 38162 31320 40000 31376
rect 38101 31318 40000 31320
rect 38101 31315 38167 31318
rect 39200 31228 40000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 38101 30698 38167 30701
rect 39200 30698 40000 30788
rect 38101 30696 40000 30698
rect 38101 30640 38106 30696
rect 38162 30640 40000 30696
rect 38101 30638 40000 30640
rect 38101 30635 38167 30638
rect 11881 30562 11947 30565
rect 16757 30562 16823 30565
rect 11881 30560 16823 30562
rect 11881 30504 11886 30560
rect 11942 30504 16762 30560
rect 16818 30504 16823 30560
rect 39200 30548 40000 30638
rect 11881 30502 16823 30504
rect 11881 30499 11947 30502
rect 16757 30499 16823 30502
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 30741 30426 30807 30429
rect 31518 30426 31524 30428
rect 30741 30424 31524 30426
rect 30741 30368 30746 30424
rect 30802 30368 31524 30424
rect 30741 30366 31524 30368
rect 30741 30363 30807 30366
rect 31518 30364 31524 30366
rect 31588 30364 31594 30428
rect 27245 30290 27311 30293
rect 27705 30290 27771 30293
rect 27245 30288 27771 30290
rect 27245 30232 27250 30288
rect 27306 30232 27710 30288
rect 27766 30232 27771 30288
rect 27245 30230 27771 30232
rect 27245 30227 27311 30230
rect 27705 30227 27771 30230
rect 0 29868 800 30108
rect 38101 30018 38167 30021
rect 39200 30018 40000 30108
rect 38101 30016 40000 30018
rect 38101 29960 38106 30016
rect 38162 29960 40000 30016
rect 38101 29958 40000 29960
rect 38101 29955 38167 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 26969 29882 27035 29885
rect 28073 29882 28139 29885
rect 26969 29880 28139 29882
rect 26969 29824 26974 29880
rect 27030 29824 28078 29880
rect 28134 29824 28139 29880
rect 39200 29868 40000 29958
rect 26969 29822 28139 29824
rect 26969 29819 27035 29822
rect 28073 29819 28139 29822
rect 12249 29474 12315 29477
rect 13629 29474 13695 29477
rect 12249 29472 13695 29474
rect 0 29188 800 29428
rect 12249 29416 12254 29472
rect 12310 29416 13634 29472
rect 13690 29416 13695 29472
rect 12249 29414 13695 29416
rect 12249 29411 12315 29414
rect 13629 29411 13695 29414
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 25497 29338 25563 29341
rect 28441 29338 28507 29341
rect 25497 29336 28507 29338
rect 25497 29280 25502 29336
rect 25558 29280 28446 29336
rect 28502 29280 28507 29336
rect 25497 29278 28507 29280
rect 25497 29275 25563 29278
rect 28441 29275 28507 29278
rect 37181 29338 37247 29341
rect 39200 29338 40000 29428
rect 37181 29336 40000 29338
rect 37181 29280 37186 29336
rect 37242 29280 40000 29336
rect 37181 29278 40000 29280
rect 37181 29275 37247 29278
rect 37549 29202 37615 29205
rect 12390 29200 37615 29202
rect 12390 29144 37554 29200
rect 37610 29144 37615 29200
rect 39200 29188 40000 29278
rect 12390 29142 37615 29144
rect 4153 29066 4219 29069
rect 5441 29066 5507 29069
rect 12390 29066 12450 29142
rect 37549 29139 37615 29142
rect 4153 29064 12450 29066
rect 4153 29008 4158 29064
rect 4214 29008 5446 29064
rect 5502 29008 12450 29064
rect 4153 29006 12450 29008
rect 26049 29066 26115 29069
rect 30373 29066 30439 29069
rect 26049 29064 30439 29066
rect 26049 29008 26054 29064
rect 26110 29008 30378 29064
rect 30434 29008 30439 29064
rect 26049 29006 30439 29008
rect 4153 29003 4219 29006
rect 5441 29003 5507 29006
rect 26049 29003 26115 29006
rect 30373 29003 30439 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28508 800 28748
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 39200 27828 40000 28068
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 27337 27570 27403 27573
rect 28165 27570 28231 27573
rect 27337 27568 28231 27570
rect 27337 27512 27342 27568
rect 27398 27512 28170 27568
rect 28226 27512 28231 27568
rect 27337 27510 28231 27512
rect 27337 27507 27403 27510
rect 28165 27507 28231 27510
rect 26325 27434 26391 27437
rect 27889 27434 27955 27437
rect 26325 27432 27955 27434
rect 26325 27376 26330 27432
rect 26386 27376 27894 27432
rect 27950 27376 27955 27432
rect 26325 27374 27955 27376
rect 26325 27371 26391 27374
rect 27889 27371 27955 27374
rect 27429 27298 27495 27301
rect 28349 27298 28415 27301
rect 27429 27296 28415 27298
rect 27429 27240 27434 27296
rect 27490 27240 28354 27296
rect 28410 27240 28415 27296
rect 27429 27238 28415 27240
rect 27429 27235 27495 27238
rect 28349 27235 28415 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 39200 27148 40000 27388
rect 23565 26890 23631 26893
rect 36261 26890 36327 26893
rect 23565 26888 36327 26890
rect 23565 26832 23570 26888
rect 23626 26832 36266 26888
rect 36322 26832 36327 26888
rect 23565 26830 36327 26832
rect 23565 26827 23631 26830
rect 36261 26827 36327 26830
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 39200 26468 40000 26708
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25938 800 26028
rect 2865 25938 2931 25941
rect 0 25936 2931 25938
rect 0 25880 2870 25936
rect 2926 25880 2931 25936
rect 0 25878 2931 25880
rect 0 25788 800 25878
rect 2865 25875 2931 25878
rect 38101 25938 38167 25941
rect 39200 25938 40000 26028
rect 38101 25936 40000 25938
rect 38101 25880 38106 25936
rect 38162 25880 40000 25936
rect 38101 25878 40000 25880
rect 38101 25875 38167 25878
rect 39200 25788 40000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25108 800 25348
rect 2313 25258 2379 25261
rect 21265 25258 21331 25261
rect 21766 25258 21772 25260
rect 2313 25256 21772 25258
rect 2313 25200 2318 25256
rect 2374 25200 21270 25256
rect 21326 25200 21772 25256
rect 2313 25198 21772 25200
rect 2313 25195 2379 25198
rect 21265 25195 21331 25198
rect 21766 25196 21772 25198
rect 21836 25196 21842 25260
rect 39200 25108 40000 25348
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 39200 24428 40000 24668
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 38101 23898 38167 23901
rect 39200 23898 40000 23988
rect 38101 23896 40000 23898
rect 38101 23840 38106 23896
rect 38162 23840 40000 23896
rect 38101 23838 40000 23840
rect 38101 23835 38167 23838
rect 39200 23748 40000 23838
rect 14365 23490 14431 23493
rect 20662 23490 20668 23492
rect 14365 23488 20668 23490
rect 14365 23432 14370 23488
rect 14426 23432 20668 23488
rect 14365 23430 20668 23432
rect 14365 23427 14431 23430
rect 20662 23428 20668 23430
rect 20732 23428 20738 23492
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23068 800 23308
rect 21173 23218 21239 23221
rect 28441 23218 28507 23221
rect 21173 23216 28507 23218
rect 21173 23160 21178 23216
rect 21234 23160 28446 23216
rect 28502 23160 28507 23216
rect 21173 23158 28507 23160
rect 21173 23155 21239 23158
rect 28441 23155 28507 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 20529 22538 20595 22541
rect 35985 22538 36051 22541
rect 20529 22536 36051 22538
rect 20529 22480 20534 22536
rect 20590 22480 35990 22536
rect 36046 22480 36051 22536
rect 20529 22478 36051 22480
rect 20529 22475 20595 22478
rect 35985 22475 36051 22478
rect 36721 22538 36787 22541
rect 39200 22538 40000 22628
rect 36721 22536 40000 22538
rect 36721 22480 36726 22536
rect 36782 22480 40000 22536
rect 36721 22478 40000 22480
rect 36721 22475 36787 22478
rect 23013 22404 23079 22405
rect 23013 22400 23060 22404
rect 23124 22402 23130 22404
rect 23013 22344 23018 22400
rect 23013 22340 23060 22344
rect 23124 22342 23170 22402
rect 39200 22388 40000 22478
rect 23124 22340 23130 22342
rect 23013 22339 23079 22340
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 21449 22266 21515 22269
rect 21449 22264 23674 22266
rect 21449 22208 21454 22264
rect 21510 22208 23674 22264
rect 21449 22206 23674 22208
rect 21449 22203 21515 22206
rect 7189 22130 7255 22133
rect 7833 22130 7899 22133
rect 7189 22128 7899 22130
rect 7189 22072 7194 22128
rect 7250 22072 7838 22128
rect 7894 22072 7899 22128
rect 7189 22070 7899 22072
rect 7189 22067 7255 22070
rect 7833 22067 7899 22070
rect 10225 22130 10291 22133
rect 11329 22130 11395 22133
rect 15285 22130 15351 22133
rect 10225 22128 15351 22130
rect 10225 22072 10230 22128
rect 10286 22072 11334 22128
rect 11390 22072 15290 22128
rect 15346 22072 15351 22128
rect 10225 22070 15351 22072
rect 10225 22067 10291 22070
rect 11329 22067 11395 22070
rect 15285 22067 15351 22070
rect 23614 21994 23674 22206
rect 23933 21994 23999 21997
rect 23614 21992 23999 21994
rect 23614 21936 23938 21992
rect 23994 21936 23999 21992
rect 23614 21934 23999 21936
rect 23933 21931 23999 21934
rect 37457 21858 37523 21861
rect 39200 21858 40000 21948
rect 37457 21856 40000 21858
rect 37457 21800 37462 21856
rect 37518 21800 40000 21856
rect 37457 21798 40000 21800
rect 37457 21795 37523 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 39200 21708 40000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 38101 21178 38167 21181
rect 39200 21178 40000 21268
rect 38101 21176 40000 21178
rect 38101 21120 38106 21176
rect 38162 21120 40000 21176
rect 38101 21118 40000 21120
rect 38101 21115 38167 21118
rect 39200 21028 40000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 13629 20498 13695 20501
rect 17861 20498 17927 20501
rect 13629 20496 17927 20498
rect 13629 20440 13634 20496
rect 13690 20440 17866 20496
rect 17922 20440 17927 20496
rect 13629 20438 17927 20440
rect 13629 20435 13695 20438
rect 17861 20435 17927 20438
rect 27429 20498 27495 20501
rect 28257 20498 28323 20501
rect 27429 20496 28323 20498
rect 27429 20440 27434 20496
rect 27490 20440 28262 20496
rect 28318 20440 28323 20496
rect 27429 20438 28323 20440
rect 27429 20435 27495 20438
rect 28257 20435 28323 20438
rect 37089 20498 37155 20501
rect 39200 20498 40000 20588
rect 37089 20496 40000 20498
rect 37089 20440 37094 20496
rect 37150 20440 40000 20496
rect 37089 20438 40000 20440
rect 37089 20435 37155 20438
rect 25129 20362 25195 20365
rect 26141 20362 26207 20365
rect 27889 20362 27955 20365
rect 25129 20360 27955 20362
rect 25129 20304 25134 20360
rect 25190 20304 26146 20360
rect 26202 20304 27894 20360
rect 27950 20304 27955 20360
rect 25129 20302 27955 20304
rect 25129 20299 25195 20302
rect 26141 20299 26207 20302
rect 27889 20299 27955 20302
rect 28257 20362 28323 20365
rect 28901 20362 28967 20365
rect 28257 20360 28967 20362
rect 28257 20304 28262 20360
rect 28318 20304 28906 20360
rect 28962 20304 28967 20360
rect 28257 20302 28967 20304
rect 28257 20299 28323 20302
rect 28901 20299 28967 20302
rect 31293 20362 31359 20365
rect 31518 20362 31524 20364
rect 31293 20360 31524 20362
rect 31293 20304 31298 20360
rect 31354 20304 31524 20360
rect 31293 20302 31524 20304
rect 31293 20299 31359 20302
rect 31518 20300 31524 20302
rect 31588 20300 31594 20364
rect 39200 20348 40000 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 20713 20092 20779 20093
rect 20662 20028 20668 20092
rect 20732 20090 20779 20092
rect 20732 20088 20824 20090
rect 20774 20032 20824 20088
rect 20732 20030 20824 20032
rect 20732 20028 20779 20030
rect 20713 20027 20779 20028
rect 22369 19954 22435 19957
rect 28901 19954 28967 19957
rect 22369 19952 28967 19954
rect 0 19818 800 19908
rect 22369 19896 22374 19952
rect 22430 19896 28906 19952
rect 28962 19896 28967 19952
rect 22369 19894 28967 19896
rect 22369 19891 22435 19894
rect 28901 19891 28967 19894
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19668 800 19758
rect 1853 19755 1919 19758
rect 15101 19818 15167 19821
rect 17309 19818 17375 19821
rect 15101 19816 17375 19818
rect 15101 19760 15106 19816
rect 15162 19760 17314 19816
rect 17370 19760 17375 19816
rect 15101 19758 17375 19760
rect 15101 19755 15167 19758
rect 17309 19755 17375 19758
rect 20713 19818 20779 19821
rect 31477 19818 31543 19821
rect 20713 19816 31543 19818
rect 20713 19760 20718 19816
rect 20774 19760 31482 19816
rect 31538 19760 31543 19816
rect 20713 19758 31543 19760
rect 20713 19755 20779 19758
rect 31477 19755 31543 19758
rect 39200 19668 40000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 11881 19546 11947 19549
rect 15009 19546 15075 19549
rect 11881 19544 15075 19546
rect 11881 19488 11886 19544
rect 11942 19488 15014 19544
rect 15070 19488 15075 19544
rect 11881 19486 15075 19488
rect 11881 19483 11947 19486
rect 15009 19483 15075 19486
rect 16757 19546 16823 19549
rect 18597 19546 18663 19549
rect 16757 19544 18663 19546
rect 16757 19488 16762 19544
rect 16818 19488 18602 19544
rect 18658 19488 18663 19544
rect 16757 19486 18663 19488
rect 16757 19483 16823 19486
rect 18597 19483 18663 19486
rect 13905 19410 13971 19413
rect 14365 19410 14431 19413
rect 18413 19410 18479 19413
rect 13905 19408 18479 19410
rect 13905 19352 13910 19408
rect 13966 19352 14370 19408
rect 14426 19352 18418 19408
rect 18474 19352 18479 19408
rect 13905 19350 18479 19352
rect 13905 19347 13971 19350
rect 14365 19347 14431 19350
rect 18413 19347 18479 19350
rect 0 19138 800 19228
rect 22134 19212 22140 19276
rect 22204 19274 22210 19276
rect 23013 19274 23079 19277
rect 27613 19274 27679 19277
rect 22204 19272 27679 19274
rect 22204 19216 23018 19272
rect 23074 19216 27618 19272
rect 27674 19216 27679 19272
rect 22204 19214 27679 19216
rect 22204 19212 22210 19214
rect 23013 19211 23079 19214
rect 27613 19211 27679 19214
rect 34973 19274 35039 19277
rect 35382 19274 35388 19276
rect 34973 19272 35388 19274
rect 34973 19216 34978 19272
rect 35034 19216 35388 19272
rect 34973 19214 35388 19216
rect 34973 19211 35039 19214
rect 35382 19212 35388 19214
rect 35452 19212 35458 19276
rect 2129 19138 2195 19141
rect 0 19136 2195 19138
rect 0 19080 2134 19136
rect 2190 19080 2195 19136
rect 0 19078 2195 19080
rect 0 18988 800 19078
rect 2129 19075 2195 19078
rect 35433 19138 35499 19141
rect 39200 19138 40000 19228
rect 35433 19136 40000 19138
rect 35433 19080 35438 19136
rect 35494 19080 40000 19136
rect 35433 19078 40000 19080
rect 35433 19075 35499 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 39200 18988 40000 19078
rect 30005 18866 30071 18869
rect 32029 18866 32095 18869
rect 30005 18864 32095 18866
rect 30005 18808 30010 18864
rect 30066 18808 32034 18864
rect 32090 18808 32095 18864
rect 30005 18806 32095 18808
rect 30005 18803 30071 18806
rect 32029 18803 32095 18806
rect 34513 18730 34579 18733
rect 34881 18730 34947 18733
rect 34513 18728 34947 18730
rect 34513 18672 34518 18728
rect 34574 18672 34886 18728
rect 34942 18672 34947 18728
rect 34513 18670 34947 18672
rect 34513 18667 34579 18670
rect 34881 18667 34947 18670
rect 0 18308 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 37089 18458 37155 18461
rect 39200 18458 40000 18548
rect 37089 18456 40000 18458
rect 37089 18400 37094 18456
rect 37150 18400 40000 18456
rect 37089 18398 40000 18400
rect 37089 18395 37155 18398
rect 39200 18308 40000 18398
rect 27245 18050 27311 18053
rect 33225 18050 33291 18053
rect 27245 18048 33291 18050
rect 27245 17992 27250 18048
rect 27306 17992 33230 18048
rect 33286 17992 33291 18048
rect 27245 17990 33291 17992
rect 27245 17987 27311 17990
rect 33225 17987 33291 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17628 800 17718
rect 2773 17715 2839 17718
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 16948 800 17188
rect 36721 17098 36787 17101
rect 39200 17098 40000 17188
rect 36721 17096 40000 17098
rect 36721 17040 36726 17096
rect 36782 17040 40000 17096
rect 36721 17038 40000 17040
rect 36721 17035 36787 17038
rect 39200 16948 40000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19241 16690 19307 16693
rect 23054 16690 23060 16692
rect 19241 16688 23060 16690
rect 19241 16632 19246 16688
rect 19302 16632 23060 16688
rect 19241 16630 23060 16632
rect 19241 16627 19307 16630
rect 23054 16628 23060 16630
rect 23124 16628 23130 16692
rect 27245 16690 27311 16693
rect 28625 16690 28691 16693
rect 27245 16688 28691 16690
rect 27245 16632 27250 16688
rect 27306 16632 28630 16688
rect 28686 16632 28691 16688
rect 27245 16630 28691 16632
rect 27245 16627 27311 16630
rect 28625 16627 28691 16630
rect 23197 16554 23263 16557
rect 31937 16554 32003 16557
rect 23197 16552 32003 16554
rect 23197 16496 23202 16552
rect 23258 16496 31942 16552
rect 31998 16496 32003 16552
rect 23197 16494 32003 16496
rect 23197 16491 23263 16494
rect 31937 16491 32003 16494
rect 38101 16418 38167 16421
rect 39200 16418 40000 16508
rect 38101 16416 40000 16418
rect 38101 16360 38106 16416
rect 38162 16360 40000 16416
rect 38101 16358 40000 16360
rect 38101 16355 38167 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 39200 16268 40000 16358
rect 24209 16146 24275 16149
rect 24710 16146 24716 16148
rect 24209 16144 24716 16146
rect 24209 16088 24214 16144
rect 24270 16088 24716 16144
rect 24209 16086 24716 16088
rect 24209 16083 24275 16086
rect 24710 16084 24716 16086
rect 24780 16146 24786 16148
rect 27061 16146 27127 16149
rect 24780 16144 27127 16146
rect 24780 16088 27066 16144
rect 27122 16088 27127 16144
rect 24780 16086 27127 16088
rect 24780 16084 24786 16086
rect 27061 16083 27127 16086
rect 0 15738 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15588 800 15678
rect 1393 15675 1459 15678
rect 35249 15602 35315 15605
rect 35382 15602 35388 15604
rect 35249 15600 35388 15602
rect 35249 15544 35254 15600
rect 35310 15544 35388 15600
rect 35249 15542 35388 15544
rect 35249 15539 35315 15542
rect 35382 15540 35388 15542
rect 35452 15540 35458 15604
rect 39200 15588 40000 15828
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 14908 800 15148
rect 38101 15058 38167 15061
rect 39200 15058 40000 15148
rect 38101 15056 40000 15058
rect 38101 15000 38106 15056
rect 38162 15000 40000 15056
rect 38101 14998 40000 15000
rect 38101 14995 38167 14998
rect 39200 14908 40000 14998
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 20897 14650 20963 14653
rect 22134 14650 22140 14652
rect 20897 14648 22140 14650
rect 20897 14592 20902 14648
rect 20958 14592 22140 14648
rect 20897 14590 22140 14592
rect 20897 14587 20963 14590
rect 22134 14588 22140 14590
rect 22204 14588 22210 14652
rect 0 14378 800 14468
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14228 800 14318
rect 1393 14315 1459 14318
rect 37089 14378 37155 14381
rect 39200 14378 40000 14468
rect 37089 14376 40000 14378
rect 37089 14320 37094 14376
rect 37150 14320 40000 14376
rect 37089 14318 40000 14320
rect 37089 14315 37155 14318
rect 39200 14228 40000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 34462 13772 34468 13836
rect 34532 13834 34538 13836
rect 35157 13834 35223 13837
rect 34532 13832 35223 13834
rect 34532 13776 35162 13832
rect 35218 13776 35223 13832
rect 34532 13774 35223 13776
rect 34532 13772 34538 13774
rect 35157 13771 35223 13774
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13548 800 13638
rect 2773 13635 2839 13638
rect 38101 13698 38167 13701
rect 39200 13698 40000 13788
rect 38101 13696 40000 13698
rect 38101 13640 38106 13696
rect 38162 13640 40000 13696
rect 38101 13638 40000 13640
rect 38101 13635 38167 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 39200 13548 40000 13638
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 30281 12882 30347 12885
rect 32397 12882 32463 12885
rect 30281 12880 32463 12882
rect 30281 12824 30286 12880
rect 30342 12824 32402 12880
rect 32458 12824 32463 12880
rect 39200 12868 40000 13108
rect 30281 12822 32463 12824
rect 30281 12819 30347 12822
rect 32397 12819 32463 12822
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 19057 12474 19123 12477
rect 19057 12472 23674 12474
rect 0 12338 800 12428
rect 19057 12416 19062 12472
rect 19118 12416 23674 12472
rect 19057 12414 23674 12416
rect 19057 12411 19123 12414
rect 23614 12341 23674 12414
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 23614 12338 23723 12341
rect 27337 12338 27403 12341
rect 32489 12338 32555 12341
rect 23614 12336 32555 12338
rect 23614 12280 23662 12336
rect 23718 12280 27342 12336
rect 27398 12280 32494 12336
rect 32550 12280 32555 12336
rect 23614 12278 32555 12280
rect 0 12188 800 12278
rect 2773 12275 2839 12278
rect 23657 12275 23723 12278
rect 27337 12275 27403 12278
rect 32489 12275 32555 12278
rect 30465 12202 30531 12205
rect 34462 12202 34468 12204
rect 30465 12200 34468 12202
rect 30465 12144 30470 12200
rect 30526 12144 34468 12200
rect 30465 12142 34468 12144
rect 30465 12139 30531 12142
rect 34462 12140 34468 12142
rect 34532 12140 34538 12204
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11658 800 11748
rect 30966 11732 30972 11796
rect 31036 11794 31042 11796
rect 36721 11794 36787 11797
rect 31036 11792 36787 11794
rect 31036 11736 36726 11792
rect 36782 11736 36787 11792
rect 31036 11734 36787 11736
rect 31036 11732 31042 11734
rect 36721 11731 36787 11734
rect 2037 11658 2103 11661
rect 0 11656 2103 11658
rect 0 11600 2042 11656
rect 2098 11600 2103 11656
rect 0 11598 2103 11600
rect 0 11508 800 11598
rect 2037 11595 2103 11598
rect 38101 11658 38167 11661
rect 39200 11658 40000 11748
rect 38101 11656 40000 11658
rect 38101 11600 38106 11656
rect 38162 11600 40000 11656
rect 38101 11598 40000 11600
rect 38101 11595 38167 11598
rect 39200 11508 40000 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 23657 11116 23723 11117
rect 23606 11052 23612 11116
rect 23676 11114 23723 11116
rect 23676 11112 23768 11114
rect 23718 11056 23768 11112
rect 23676 11054 23768 11056
rect 23676 11052 23723 11054
rect 23657 11051 23723 11052
rect 35801 10978 35867 10981
rect 39200 10978 40000 11068
rect 35801 10976 40000 10978
rect 35801 10920 35806 10976
rect 35862 10920 40000 10976
rect 35801 10918 40000 10920
rect 35801 10915 35867 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 21541 10842 21607 10845
rect 24117 10842 24183 10845
rect 21541 10840 24183 10842
rect 21541 10784 21546 10840
rect 21602 10784 24122 10840
rect 24178 10784 24183 10840
rect 39200 10828 40000 10918
rect 21541 10782 24183 10784
rect 21541 10779 21607 10782
rect 24117 10779 24183 10782
rect 0 10148 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 38101 10298 38167 10301
rect 39200 10298 40000 10388
rect 38101 10296 40000 10298
rect 38101 10240 38106 10296
rect 38162 10240 40000 10296
rect 38101 10238 40000 10240
rect 38101 10235 38167 10238
rect 39200 10148 40000 10238
rect 19333 10026 19399 10029
rect 26509 10026 26575 10029
rect 19333 10024 26575 10026
rect 19333 9968 19338 10024
rect 19394 9968 26514 10024
rect 26570 9968 26575 10024
rect 19333 9966 26575 9968
rect 19333 9963 19399 9966
rect 26509 9963 26575 9966
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 37181 9618 37247 9621
rect 39200 9618 40000 9708
rect 37181 9616 40000 9618
rect 37181 9560 37186 9616
rect 37242 9560 40000 9616
rect 37181 9558 40000 9560
rect 37181 9555 37247 9558
rect 39200 9468 40000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 9028
rect 1853 8938 1919 8941
rect 0 8936 1919 8938
rect 0 8880 1858 8936
rect 1914 8880 1919 8936
rect 0 8878 1919 8880
rect 0 8788 800 8878
rect 1853 8875 1919 8878
rect 20069 8938 20135 8941
rect 20253 8938 20319 8941
rect 22277 8938 22343 8941
rect 20069 8936 22343 8938
rect 20069 8880 20074 8936
rect 20130 8880 20258 8936
rect 20314 8880 22282 8936
rect 22338 8880 22343 8936
rect 20069 8878 22343 8880
rect 20069 8875 20135 8878
rect 20253 8875 20319 8878
rect 22277 8875 22343 8878
rect 24761 8938 24827 8941
rect 26141 8938 26207 8941
rect 24761 8936 26207 8938
rect 24761 8880 24766 8936
rect 24822 8880 26146 8936
rect 26202 8880 26207 8936
rect 24761 8878 26207 8880
rect 24761 8875 24827 8878
rect 26141 8875 26207 8878
rect 25589 8802 25655 8805
rect 27981 8802 28047 8805
rect 25589 8800 28047 8802
rect 25589 8744 25594 8800
rect 25650 8744 27986 8800
rect 28042 8744 28047 8800
rect 39200 8788 40000 9028
rect 25589 8742 28047 8744
rect 25589 8739 25655 8742
rect 27981 8739 28047 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8258 800 8348
rect 3969 8258 4035 8261
rect 0 8256 4035 8258
rect 0 8200 3974 8256
rect 4030 8200 4035 8256
rect 0 8198 4035 8200
rect 0 8108 800 8198
rect 3969 8195 4035 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 39200 8108 40000 8348
rect 21449 7986 21515 7989
rect 27797 7986 27863 7989
rect 21449 7984 27863 7986
rect 21449 7928 21454 7984
rect 21510 7928 27802 7984
rect 27858 7928 27863 7984
rect 21449 7926 27863 7928
rect 21449 7923 21515 7926
rect 27797 7923 27863 7926
rect 21081 7850 21147 7853
rect 27153 7850 27219 7853
rect 21081 7848 27219 7850
rect 21081 7792 21086 7848
rect 21142 7792 27158 7848
rect 27214 7792 27219 7848
rect 21081 7790 27219 7792
rect 21081 7787 21147 7790
rect 27153 7787 27219 7790
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 2773 7578 2839 7581
rect 0 7576 2839 7578
rect 0 7520 2778 7576
rect 2834 7520 2839 7576
rect 0 7518 2839 7520
rect 0 7428 800 7518
rect 2773 7515 2839 7518
rect 20897 7578 20963 7581
rect 23606 7578 23612 7580
rect 20897 7576 23612 7578
rect 20897 7520 20902 7576
rect 20958 7520 23612 7576
rect 20897 7518 23612 7520
rect 20897 7515 20963 7518
rect 23606 7516 23612 7518
rect 23676 7516 23682 7580
rect 24710 7380 24716 7444
rect 24780 7442 24786 7444
rect 27429 7442 27495 7445
rect 24780 7440 27495 7442
rect 24780 7384 27434 7440
rect 27490 7384 27495 7440
rect 39200 7428 40000 7668
rect 24780 7382 27495 7384
rect 24780 7380 24786 7382
rect 27429 7379 27495 7382
rect 19425 7306 19491 7309
rect 23657 7306 23723 7309
rect 24209 7306 24275 7309
rect 19425 7304 24275 7306
rect 19425 7248 19430 7304
rect 19486 7248 23662 7304
rect 23718 7248 24214 7304
rect 24270 7248 24275 7304
rect 19425 7246 24275 7248
rect 19425 7243 19491 7246
rect 23657 7243 23723 7246
rect 24209 7243 24275 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6748 800 6988
rect 22134 6972 22140 7036
rect 22204 7034 22210 7036
rect 26325 7034 26391 7037
rect 22204 7032 26391 7034
rect 22204 6976 26330 7032
rect 26386 6976 26391 7032
rect 22204 6974 26391 6976
rect 22204 6972 22210 6974
rect 26325 6971 26391 6974
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6218 800 6308
rect 2773 6218 2839 6221
rect 0 6216 2839 6218
rect 0 6160 2778 6216
rect 2834 6160 2839 6216
rect 0 6158 2839 6160
rect 0 6068 800 6158
rect 2773 6155 2839 6158
rect 38009 6218 38075 6221
rect 39200 6218 40000 6308
rect 38009 6216 40000 6218
rect 38009 6160 38014 6216
rect 38070 6160 40000 6216
rect 38009 6158 40000 6160
rect 38009 6155 38075 6158
rect 39200 6068 40000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 37181 5538 37247 5541
rect 39200 5538 40000 5628
rect 37181 5536 40000 5538
rect 37181 5480 37186 5536
rect 37242 5480 40000 5536
rect 37181 5478 40000 5480
rect 37181 5475 37247 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 39200 5388 40000 5478
rect 21214 5204 21220 5268
rect 21284 5266 21290 5268
rect 36629 5266 36695 5269
rect 21284 5264 36695 5266
rect 21284 5208 36634 5264
rect 36690 5208 36695 5264
rect 21284 5206 36695 5208
rect 21284 5204 21290 5206
rect 36629 5203 36695 5206
rect 0 4858 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 1761 4858 1827 4861
rect 0 4856 1827 4858
rect 0 4800 1766 4856
rect 1822 4800 1827 4856
rect 0 4798 1827 4800
rect 0 4708 800 4798
rect 1761 4795 1827 4798
rect 39200 4708 40000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4268
rect 3417 4178 3483 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4028 800 4118
rect 3417 4115 3483 4118
rect 37549 4178 37615 4181
rect 39200 4178 40000 4268
rect 37549 4176 40000 4178
rect 37549 4120 37554 4176
rect 37610 4120 40000 4176
rect 37549 4118 40000 4120
rect 37549 4115 37615 4118
rect 5165 4042 5231 4045
rect 7230 4042 7236 4044
rect 5165 4040 7236 4042
rect 5165 3984 5170 4040
rect 5226 3984 7236 4040
rect 5165 3982 7236 3984
rect 5165 3979 5231 3982
rect 7230 3980 7236 3982
rect 7300 3980 7306 4044
rect 20713 4042 20779 4045
rect 20846 4042 20852 4044
rect 20713 4040 20852 4042
rect 20713 3984 20718 4040
rect 20774 3984 20852 4040
rect 20713 3982 20852 3984
rect 20713 3979 20779 3982
rect 20846 3980 20852 3982
rect 20916 3980 20922 4044
rect 21766 3980 21772 4044
rect 21836 4042 21842 4044
rect 24669 4042 24735 4045
rect 21836 4040 24735 4042
rect 21836 3984 24674 4040
rect 24730 3984 24735 4040
rect 39200 4028 40000 4118
rect 21836 3982 24735 3984
rect 21836 3980 21842 3982
rect 24669 3979 24735 3982
rect 23054 3844 23060 3908
rect 23124 3906 23130 3908
rect 31385 3906 31451 3909
rect 23124 3904 31451 3906
rect 23124 3848 31390 3904
rect 31446 3848 31451 3904
rect 23124 3846 31451 3848
rect 23124 3844 23130 3846
rect 31385 3843 31451 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 39200 3348 40000 3588
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 0 2818 800 2908
rect 2773 2818 2839 2821
rect 0 2816 2839 2818
rect 0 2760 2778 2816
rect 2834 2760 2839 2816
rect 0 2758 2839 2760
rect 0 2668 800 2758
rect 2773 2755 2839 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 39200 2668 40000 2908
rect 0 2138 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 1393 2138 1459 2141
rect 0 2136 1459 2138
rect 0 2080 1398 2136
rect 1454 2080 1459 2136
rect 0 2078 1459 2080
rect 0 1988 800 2078
rect 1393 2075 1459 2078
rect 35801 2138 35867 2141
rect 39200 2138 40000 2228
rect 35801 2136 40000 2138
rect 35801 2080 35806 2136
rect 35862 2080 40000 2136
rect 35801 2078 40000 2080
rect 35801 2075 35867 2078
rect 39200 1988 40000 2078
rect 0 1458 800 1548
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1308 800 1398
rect 2865 1395 2931 1398
rect 0 628 800 868
rect 37089 778 37155 781
rect 39200 778 40000 868
rect 37089 776 40000 778
rect 37089 720 37094 776
rect 37150 720 40000 776
rect 37089 718 40000 720
rect 37089 715 37155 718
rect 39200 628 40000 718
rect 35157 98 35223 101
rect 39200 98 40000 188
rect 35157 96 40000 98
rect 35157 40 35162 96
rect 35218 40 40000 96
rect 35157 38 40000 40
rect 35157 35 35223 38
rect 39200 -52 40000 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 7236 36816 7300 36820
rect 7236 36760 7250 36816
rect 7250 36760 7300 36816
rect 7236 36756 7300 36760
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 30972 35940 31036 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 21220 35532 21284 35596
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 20852 32948 20916 33012
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 31524 30364 31588 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 21772 25196 21836 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 20668 23428 20732 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 23060 22400 23124 22404
rect 23060 22344 23074 22400
rect 23074 22344 23124 22400
rect 23060 22340 23124 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 31524 20300 31588 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 20668 20088 20732 20092
rect 20668 20032 20718 20088
rect 20718 20032 20732 20088
rect 20668 20028 20732 20032
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 22140 19212 22204 19276
rect 35388 19212 35452 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 23060 16628 23124 16692
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 24716 16084 24780 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 35388 15540 35452 15604
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 22140 14588 22204 14652
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 34468 13772 34532 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 34468 12140 34532 12204
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 30972 11732 31036 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 23612 11112 23676 11116
rect 23612 11056 23662 11112
rect 23662 11056 23676 11112
rect 23612 11052 23676 11056
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 23612 7516 23676 7580
rect 24716 7380 24780 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 22140 6972 22204 7036
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 21220 5204 21284 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 7236 3980 7300 4044
rect 20852 3980 20916 4044
rect 21772 3980 21836 4044
rect 23060 3844 23124 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 7235 36820 7301 36821
rect 7235 36756 7236 36820
rect 7300 36756 7301 36820
rect 7235 36755 7301 36756
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 7238 4045 7298 36755
rect 19568 35936 19888 36960
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 30971 36004 31037 36005
rect 30971 35940 30972 36004
rect 31036 35940 31037 36004
rect 30971 35939 31037 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 21219 35596 21285 35597
rect 21219 35532 21220 35596
rect 21284 35532 21285 35596
rect 21219 35531 21285 35532
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 20851 33012 20917 33013
rect 20851 32948 20852 33012
rect 20916 32948 20917 33012
rect 20851 32947 20917 32948
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 20667 23492 20733 23493
rect 20667 23428 20668 23492
rect 20732 23428 20733 23492
rect 20667 23427 20733 23428
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 20670 20093 20730 23427
rect 20667 20092 20733 20093
rect 20667 20028 20668 20092
rect 20732 20028 20733 20092
rect 20667 20027 20733 20028
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 7235 4044 7301 4045
rect 7235 3980 7236 4044
rect 7300 3980 7301 4044
rect 7235 3979 7301 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 20854 4045 20914 32947
rect 21222 5269 21282 35531
rect 21771 25260 21837 25261
rect 21771 25196 21772 25260
rect 21836 25196 21837 25260
rect 21771 25195 21837 25196
rect 21219 5268 21285 5269
rect 21219 5204 21220 5268
rect 21284 5204 21285 5268
rect 21219 5203 21285 5204
rect 21774 4045 21834 25195
rect 23059 22404 23125 22405
rect 23059 22340 23060 22404
rect 23124 22340 23125 22404
rect 23059 22339 23125 22340
rect 22139 19276 22205 19277
rect 22139 19212 22140 19276
rect 22204 19212 22205 19276
rect 22139 19211 22205 19212
rect 22142 14653 22202 19211
rect 23062 16693 23122 22339
rect 23059 16692 23125 16693
rect 23059 16628 23060 16692
rect 23124 16628 23125 16692
rect 23059 16627 23125 16628
rect 22139 14652 22205 14653
rect 22139 14588 22140 14652
rect 22204 14588 22205 14652
rect 22139 14587 22205 14588
rect 22142 7037 22202 14587
rect 22139 7036 22205 7037
rect 22139 6972 22140 7036
rect 22204 6972 22205 7036
rect 22139 6971 22205 6972
rect 20851 4044 20917 4045
rect 20851 3980 20852 4044
rect 20916 3980 20917 4044
rect 20851 3979 20917 3980
rect 21771 4044 21837 4045
rect 21771 3980 21772 4044
rect 21836 3980 21837 4044
rect 21771 3979 21837 3980
rect 23062 3909 23122 16627
rect 24715 16148 24781 16149
rect 24715 16084 24716 16148
rect 24780 16084 24781 16148
rect 24715 16083 24781 16084
rect 23611 11116 23677 11117
rect 23611 11052 23612 11116
rect 23676 11052 23677 11116
rect 23611 11051 23677 11052
rect 23614 7581 23674 11051
rect 23611 7580 23677 7581
rect 23611 7516 23612 7580
rect 23676 7516 23677 7580
rect 23611 7515 23677 7516
rect 24718 7445 24778 16083
rect 30974 11797 31034 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 31523 30428 31589 30429
rect 31523 30364 31524 30428
rect 31588 30364 31589 30428
rect 31523 30363 31589 30364
rect 31526 20365 31586 30363
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 31523 20364 31589 20365
rect 31523 20300 31524 20364
rect 31588 20300 31589 20364
rect 31523 20299 31589 20300
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 35387 19276 35453 19277
rect 35387 19212 35388 19276
rect 35452 19212 35453 19276
rect 35387 19211 35453 19212
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 35390 15605 35450 19211
rect 35387 15604 35453 15605
rect 35387 15540 35388 15604
rect 35452 15540 35453 15604
rect 35387 15539 35453 15540
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34467 13836 34533 13837
rect 34467 13772 34468 13836
rect 34532 13772 34533 13836
rect 34467 13771 34533 13772
rect 34470 12205 34530 13771
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34467 12204 34533 12205
rect 34467 12140 34468 12204
rect 34532 12140 34533 12204
rect 34467 12139 34533 12140
rect 30971 11796 31037 11797
rect 30971 11732 30972 11796
rect 31036 11732 31037 11796
rect 30971 11731 31037 11732
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 24715 7444 24781 7445
rect 24715 7380 24716 7444
rect 24780 7380 24781 7444
rect 24715 7379 24781 7380
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 23059 3908 23125 3909
rect 23059 3844 23060 3908
rect 23124 3844 23125 3908
rect 23059 3843 23125 3844
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1644511149
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1644511149
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_172
timestamp 1644511149
transform 1 0 16928 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_188 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1644511149
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1644511149
transform 1 0 22080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_235
timestamp 1644511149
transform 1 0 22724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_242 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_259
timestamp 1644511149
transform 1 0 24932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 1644511149
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1644511149
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_48
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1644511149
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_246
timestamp 1644511149
transform 1 0 23736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1644511149
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_321
timestamp 1644511149
transform 1 0 30636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1644511149
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_358
timestamp 1644511149
transform 1 0 34040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_366
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_60
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1644511149
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_131
timestamp 1644511149
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1644511149
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_155
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1644511149
transform 1 0 16100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_176
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_211
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1644511149
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_259
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_271
timestamp 1644511149
transform 1 0 26036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_283
timestamp 1644511149
transform 1 0 27140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_295
timestamp 1644511149
transform 1 0 28244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_317
timestamp 1644511149
transform 1 0 30268 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_346
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1644511149
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_394
timestamp 1644511149
transform 1 0 37352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_36
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_133
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_145
timestamp 1644511149
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 1644511149
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1644511149
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_207
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_258
timestamp 1644511149
transform 1 0 24840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1644511149
transform 1 0 25852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1644511149
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1644511149
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_341
timestamp 1644511149
transform 1 0 32476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_363
timestamp 1644511149
transform 1 0 34500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_396
timestamp 1644511149
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1644511149
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1644511149
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_72
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1644511149
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1644511149
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_101
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1644511149
transform 1 0 10764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1644511149
transform 1 0 11868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1644511149
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1644511149
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_174
timestamp 1644511149
transform 1 0 17112 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_180
timestamp 1644511149
transform 1 0 17664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_184
timestamp 1644511149
transform 1 0 18032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_188
timestamp 1644511149
transform 1 0 18400 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_219
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_256
timestamp 1644511149
transform 1 0 24656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1644511149
transform 1 0 26864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_292
timestamp 1644511149
transform 1 0 27968 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_337
timestamp 1644511149
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_359
timestamp 1644511149
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_372
timestamp 1644511149
transform 1 0 35328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_397
timestamp 1644511149
transform 1 0 37628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1644511149
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_35
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp 1644511149
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1644511149
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_60
timestamp 1644511149
transform 1 0 6624 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_72
timestamp 1644511149
transform 1 0 7728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1644511149
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_96
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_157
timestamp 1644511149
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1644511149
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1644511149
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1644511149
transform 1 0 22172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_242
timestamp 1644511149
transform 1 0 23368 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1644511149
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_255
timestamp 1644511149
transform 1 0 24564 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_345
timestamp 1644511149
transform 1 0 32844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_367
timestamp 1644511149
transform 1 0 34868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_371
timestamp 1644511149
transform 1 0 35236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_377
timestamp 1644511149
transform 1 0 35788 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1644511149
transform 1 0 36156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_398
timestamp 1644511149
transform 1 0 37720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1644511149
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_40
timestamp 1644511149
transform 1 0 4784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1644511149
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1644511149
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1644511149
transform 1 0 15640 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1644511149
transform 1 0 16928 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_182
timestamp 1644511149
transform 1 0 17848 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_188
timestamp 1644511149
transform 1 0 18400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_201
timestamp 1644511149
transform 1 0 19596 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_229
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_237
timestamp 1644511149
transform 1 0 22908 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1644511149
transform 1 0 24840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_272
timestamp 1644511149
transform 1 0 26128 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_284
timestamp 1644511149
transform 1 0 27232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_291
timestamp 1644511149
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1644511149
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_373
timestamp 1644511149
transform 1 0 35420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_378
timestamp 1644511149
transform 1 0 35880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_155
timestamp 1644511149
transform 1 0 15364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_176
timestamp 1644511149
transform 1 0 17296 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1644511149
transform 1 0 18308 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1644511149
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1644511149
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_215
timestamp 1644511149
transform 1 0 20884 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1644511149
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_230
timestamp 1644511149
transform 1 0 22264 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1644511149
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_251
timestamp 1644511149
transform 1 0 24196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_257
timestamp 1644511149
transform 1 0 24748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_268
timestamp 1644511149
transform 1 0 25760 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_302
timestamp 1644511149
transform 1 0 28888 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_314
timestamp 1644511149
transform 1 0 29992 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_326
timestamp 1644511149
transform 1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1644511149
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1644511149
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1644511149
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1644511149
transform 1 0 2392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1644511149
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1644511149
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_166
timestamp 1644511149
transform 1 0 16376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_176
timestamp 1644511149
transform 1 0 17296 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_184
timestamp 1644511149
transform 1 0 18032 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1644511149
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_225
timestamp 1644511149
transform 1 0 21804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_234
timestamp 1644511149
transform 1 0 22632 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1644511149
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_268
timestamp 1644511149
transform 1 0 25760 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_275
timestamp 1644511149
transform 1 0 26404 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_282
timestamp 1644511149
transform 1 0 27048 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_288
timestamp 1644511149
transform 1 0 27600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_299
timestamp 1644511149
transform 1 0 28612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_312
timestamp 1644511149
transform 1 0 29808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_324
timestamp 1644511149
transform 1 0 30912 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_336
timestamp 1644511149
transform 1 0 32016 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_348
timestamp 1644511149
transform 1 0 33120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1644511149
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_381
timestamp 1644511149
transform 1 0 36156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1644511149
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_28
timestamp 1644511149
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_40
timestamp 1644511149
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1644511149
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1644511149
transform 1 0 17572 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_188
timestamp 1644511149
transform 1 0 18400 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_194
timestamp 1644511149
transform 1 0 18952 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_201
timestamp 1644511149
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_208
timestamp 1644511149
transform 1 0 20240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1644511149
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_243
timestamp 1644511149
transform 1 0 23460 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_250
timestamp 1644511149
transform 1 0 24104 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_262
timestamp 1644511149
transform 1 0 25208 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1644511149
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_289
timestamp 1644511149
transform 1 0 27692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_315
timestamp 1644511149
transform 1 0 30084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1644511149
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_378
timestamp 1644511149
transform 1 0 35880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1644511149
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_400
timestamp 1644511149
transform 1 0 37904 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_406
timestamp 1644511149
transform 1 0 38456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_10
timestamp 1644511149
transform 1 0 2024 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1644511149
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_52
timestamp 1644511149
transform 1 0 5888 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_64
timestamp 1644511149
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1644511149
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1644511149
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_167
timestamp 1644511149
transform 1 0 16468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1644511149
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_204
timestamp 1644511149
transform 1 0 19872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_208
timestamp 1644511149
transform 1 0 20240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_219
timestamp 1644511149
transform 1 0 21252 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_227
timestamp 1644511149
transform 1 0 21988 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_239
timestamp 1644511149
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_264
timestamp 1644511149
transform 1 0 25392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_268
timestamp 1644511149
transform 1 0 25760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_276
timestamp 1644511149
transform 1 0 26496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_288
timestamp 1644511149
transform 1 0 27600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1644511149
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_312
timestamp 1644511149
transform 1 0 29808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_319
timestamp 1644511149
transform 1 0 30452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_326
timestamp 1644511149
transform 1 0 31096 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_338
timestamp 1644511149
transform 1 0 32200 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_350
timestamp 1644511149
transform 1 0 33304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1644511149
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_371
timestamp 1644511149
transform 1 0 35236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_396
timestamp 1644511149
transform 1 0 37536 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1644511149
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1644511149
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1644511149
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 1644511149
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1644511149
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_175
timestamp 1644511149
transform 1 0 17204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1644511149
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_195
timestamp 1644511149
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1644511149
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_212
timestamp 1644511149
transform 1 0 20608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_230
timestamp 1644511149
transform 1 0 22264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_234
timestamp 1644511149
transform 1 0 22632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_238
timestamp 1644511149
transform 1 0 23000 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_253
timestamp 1644511149
transform 1 0 24380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_262
timestamp 1644511149
transform 1 0 25208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_285
timestamp 1644511149
transform 1 0 27324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_296
timestamp 1644511149
transform 1 0 28336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_320
timestamp 1644511149
transform 1 0 30544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1644511149
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1644511149
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_400
timestamp 1644511149
transform 1 0 37904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1644511149
transform 1 0 38456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1644511149
transform 1 0 4048 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1644511149
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_51
timestamp 1644511149
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_63
timestamp 1644511149
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1644511149
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1644511149
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_168
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_172
timestamp 1644511149
transform 1 0 16928 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1644511149
transform 1 0 17848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 1644511149
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_201
timestamp 1644511149
transform 1 0 19596 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_210
timestamp 1644511149
transform 1 0 20424 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_225
timestamp 1644511149
transform 1 0 21804 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_236
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_244
timestamp 1644511149
transform 1 0 23552 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_260
timestamp 1644511149
transform 1 0 25024 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_268
timestamp 1644511149
transform 1 0 25760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1644511149
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_287
timestamp 1644511149
transform 1 0 27508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_315
timestamp 1644511149
transform 1 0 30084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_322
timestamp 1644511149
transform 1 0 30728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_329
timestamp 1644511149
transform 1 0 31372 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_341
timestamp 1644511149
transform 1 0 32476 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_353
timestamp 1644511149
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1644511149
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_374
timestamp 1644511149
transform 1 0 35512 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_8
timestamp 1644511149
transform 1 0 1840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_16
timestamp 1644511149
transform 1 0 2576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_20
timestamp 1644511149
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1644511149
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1644511149
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1644511149
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_189
timestamp 1644511149
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1644511149
transform 1 0 19320 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_210
timestamp 1644511149
transform 1 0 20424 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_236
timestamp 1644511149
transform 1 0 22816 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_242
timestamp 1644511149
transform 1 0 23368 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_252
timestamp 1644511149
transform 1 0 24288 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_258
timestamp 1644511149
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_265
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1644511149
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1644511149
transform 1 0 28520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_319
timestamp 1644511149
transform 1 0 30452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_326
timestamp 1644511149
transform 1 0 31096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1644511149
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_360
timestamp 1644511149
transform 1 0 34224 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_371
timestamp 1644511149
transform 1 0 35236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_378
timestamp 1644511149
transform 1 0 35880 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_384
timestamp 1644511149
transform 1 0 36432 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_398
timestamp 1644511149
transform 1 0 37720 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_406
timestamp 1644511149
transform 1 0 38456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1644511149
transform 1 0 14352 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_155
timestamp 1644511149
transform 1 0 15364 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1644511149
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 1644511149
transform 1 0 17572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1644511149
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1644511149
transform 1 0 20056 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_218
timestamp 1644511149
transform 1 0 21160 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_226
timestamp 1644511149
transform 1 0 21896 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_238
timestamp 1644511149
transform 1 0 23000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_279
timestamp 1644511149
transform 1 0 26772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_296
timestamp 1644511149
transform 1 0 28336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_313
timestamp 1644511149
transform 1 0 29900 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_326
timestamp 1644511149
transform 1 0 31096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_340
timestamp 1644511149
transform 1 0 32384 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_352
timestamp 1644511149
transform 1 0 33488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_356
timestamp 1644511149
transform 1 0 33856 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1644511149
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_370
timestamp 1644511149
transform 1 0 35144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_381
timestamp 1644511149
transform 1 0 36156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1644511149
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_8
timestamp 1644511149
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_20
timestamp 1644511149
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1644511149
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1644511149
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_143
timestamp 1644511149
transform 1 0 14260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1644511149
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1644511149
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_188
timestamp 1644511149
transform 1 0 18400 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_197
timestamp 1644511149
transform 1 0 19228 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_204
timestamp 1644511149
transform 1 0 19872 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1644511149
transform 1 0 20608 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_238
timestamp 1644511149
transform 1 0 23000 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_245
timestamp 1644511149
transform 1 0 23644 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_266
timestamp 1644511149
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1644511149
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_287
timestamp 1644511149
transform 1 0 27508 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_301
timestamp 1644511149
transform 1 0 28796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_314
timestamp 1644511149
transform 1 0 29992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_322
timestamp 1644511149
transform 1 0 30728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1644511149
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_357
timestamp 1644511149
transform 1 0 33948 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_365
timestamp 1644511149
transform 1 0 34684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1644511149
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_397
timestamp 1644511149
transform 1 0 37628 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1644511149
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_144
timestamp 1644511149
transform 1 0 14352 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_170
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1644511149
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1644511149
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_206
timestamp 1644511149
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1644511149
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_228
timestamp 1644511149
transform 1 0 22080 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_238
timestamp 1644511149
transform 1 0 23000 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_263
timestamp 1644511149
transform 1 0 25300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_274
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_281
timestamp 1644511149
transform 1 0 26956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_285
timestamp 1644511149
transform 1 0 27324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1644511149
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_312
timestamp 1644511149
transform 1 0 29808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_336
timestamp 1644511149
transform 1 0 32016 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1644511149
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_371
timestamp 1644511149
transform 1 0 35236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_378
timestamp 1644511149
transform 1 0 35880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1644511149
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_26
timestamp 1644511149
transform 1 0 3496 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_38
timestamp 1644511149
transform 1 0 4600 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1644511149
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1644511149
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1644511149
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_185
timestamp 1644511149
transform 1 0 18124 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1644511149
transform 1 0 18768 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_196
timestamp 1644511149
transform 1 0 19136 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_207
timestamp 1644511149
transform 1 0 20148 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_213
timestamp 1644511149
transform 1 0 20700 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_230
timestamp 1644511149
transform 1 0 22264 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_256
timestamp 1644511149
transform 1 0 24656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_301
timestamp 1644511149
transform 1 0 28796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_325
timestamp 1644511149
transform 1 0 31004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_342
timestamp 1644511149
transform 1 0 32568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_353
timestamp 1644511149
transform 1 0 33580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_381
timestamp 1644511149
transform 1 0 36156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1644511149
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_399
timestamp 1644511149
transform 1 0 37812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_162
timestamp 1644511149
transform 1 0 16008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_170
timestamp 1644511149
transform 1 0 16744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1644511149
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1644511149
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_204
timestamp 1644511149
transform 1 0 19872 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1644511149
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1644511149
transform 1 0 21252 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1644511149
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_262
timestamp 1644511149
transform 1 0 25208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1644511149
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1644511149
transform 1 0 26496 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_297
timestamp 1644511149
transform 1 0 28428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_312
timestamp 1644511149
transform 1 0 29808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1644511149
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_329
timestamp 1644511149
transform 1 0 31372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_342
timestamp 1644511149
transform 1 0 32568 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_356
timestamp 1644511149
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_369
timestamp 1644511149
transform 1 0 35052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_378
timestamp 1644511149
transform 1 0 35880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1644511149
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_11
timestamp 1644511149
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_23
timestamp 1644511149
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_35
timestamp 1644511149
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1644511149
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1644511149
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_158
timestamp 1644511149
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1644511149
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_182
timestamp 1644511149
transform 1 0 17848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1644511149
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_204
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_209
timestamp 1644511149
transform 1 0 20332 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_215
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_252
timestamp 1644511149
transform 1 0 24288 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_260
timestamp 1644511149
transform 1 0 25024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_269
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_285
timestamp 1644511149
transform 1 0 27324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_292
timestamp 1644511149
transform 1 0 27968 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1644511149
transform 1 0 28520 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_303
timestamp 1644511149
transform 1 0 28980 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_307
timestamp 1644511149
transform 1 0 29348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_314
timestamp 1644511149
transform 1 0 29992 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_322
timestamp 1644511149
transform 1 0 30728 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1644511149
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_342
timestamp 1644511149
transform 1 0 32568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_356
timestamp 1644511149
transform 1 0 33856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_365
timestamp 1644511149
transform 1 0 34684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_380
timestamp 1644511149
transform 1 0 36064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1644511149
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_399
timestamp 1644511149
transform 1 0 37812 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_8
timestamp 1644511149
transform 1 0 1840 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_17
timestamp 1644511149
transform 1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1644511149
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1644511149
transform 1 0 16468 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1644511149
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1644511149
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_205
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1644511149
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1644511149
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1644511149
transform 1 0 22816 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_243
timestamp 1644511149
transform 1 0 23460 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_261
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_269
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1644511149
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_284
timestamp 1644511149
transform 1 0 27232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_292
timestamp 1644511149
transform 1 0 27968 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_315
timestamp 1644511149
transform 1 0 30084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_323
timestamp 1644511149
transform 1 0 30820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_329
timestamp 1644511149
transform 1 0 31372 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_335
timestamp 1644511149
transform 1 0 31924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_346
timestamp 1644511149
transform 1 0 32936 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_352
timestamp 1644511149
transform 1 0 33488 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1644511149
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_370
timestamp 1644511149
transform 1 0 35144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_378
timestamp 1644511149
transform 1 0 35880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1644511149
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_29
timestamp 1644511149
transform 1 0 3772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_41
timestamp 1644511149
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1644511149
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_121
timestamp 1644511149
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1644511149
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1644511149
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1644511149
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_180
timestamp 1644511149
transform 1 0 17664 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1644511149
transform 1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1644511149
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_236
timestamp 1644511149
transform 1 0 22816 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_257
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_266
timestamp 1644511149
transform 1 0 25576 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_285
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_291
timestamp 1644511149
transform 1 0 27876 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_351
timestamp 1644511149
transform 1 0 33396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_362
timestamp 1644511149
transform 1 0 34408 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1644511149
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_398
timestamp 1644511149
transform 1 0 37720 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1644511149
transform 1 0 38456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1644511149
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1644511149
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1644511149
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1644511149
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1644511149
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_132
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1644511149
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_162
timestamp 1644511149
transform 1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_182
timestamp 1644511149
transform 1 0 17848 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1644511149
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_224
timestamp 1644511149
transform 1 0 21712 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_236
timestamp 1644511149
transform 1 0 22816 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_273
timestamp 1644511149
transform 1 0 26220 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_281
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_302
timestamp 1644511149
transform 1 0 28888 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_319
timestamp 1644511149
transform 1 0 30452 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_347
timestamp 1644511149
transform 1 0 33028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1644511149
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_373
timestamp 1644511149
transform 1 0 35420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_381
timestamp 1644511149
transform 1 0 36156 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_19
timestamp 1644511149
transform 1 0 2852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_26
timestamp 1644511149
transform 1 0 3496 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_38
timestamp 1644511149
transform 1 0 4600 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1644511149
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_129
timestamp 1644511149
transform 1 0 12972 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1644511149
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_143
timestamp 1644511149
transform 1 0 14260 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_147
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_154
timestamp 1644511149
transform 1 0 15272 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1644511149
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1644511149
transform 1 0 19320 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1644511149
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_242
timestamp 1644511149
transform 1 0 23368 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_254
timestamp 1644511149
transform 1 0 24472 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_294
timestamp 1644511149
transform 1 0 28152 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_302
timestamp 1644511149
transform 1 0 28888 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1644511149
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1644511149
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_322
timestamp 1644511149
transform 1 0 30728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_328
timestamp 1644511149
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_342
timestamp 1644511149
transform 1 0 32568 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_346
timestamp 1644511149
transform 1 0 32936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_367
timestamp 1644511149
transform 1 0 34868 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_377
timestamp 1644511149
transform 1 0 35788 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_398
timestamp 1644511149
transform 1 0 37720 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1644511149
transform 1 0 38456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1644511149
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_119
timestamp 1644511149
transform 1 0 12052 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_145
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_169
timestamp 1644511149
transform 1 0 16652 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_183
timestamp 1644511149
transform 1 0 17940 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_187
timestamp 1644511149
transform 1 0 18308 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1644511149
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_206
timestamp 1644511149
transform 1 0 20056 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_225
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_231
timestamp 1644511149
transform 1 0 22356 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_236
timestamp 1644511149
transform 1 0 22816 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_244
timestamp 1644511149
transform 1 0 23552 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1644511149
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_282
timestamp 1644511149
transform 1 0 27048 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_290
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_298
timestamp 1644511149
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1644511149
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_312
timestamp 1644511149
transform 1 0 29808 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_323
timestamp 1644511149
transform 1 0 30820 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_332
timestamp 1644511149
transform 1 0 31648 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1644511149
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_375
timestamp 1644511149
transform 1 0 35604 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_381
timestamp 1644511149
transform 1 0 36156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1644511149
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_12
timestamp 1644511149
transform 1 0 2208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_24
timestamp 1644511149
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_36
timestamp 1644511149
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1644511149
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1644511149
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_91
timestamp 1644511149
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_103
timestamp 1644511149
transform 1 0 10580 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_129
timestamp 1644511149
transform 1 0 12972 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_135
timestamp 1644511149
transform 1 0 13524 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_152
timestamp 1644511149
transform 1 0 15088 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_158
timestamp 1644511149
transform 1 0 15640 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1644511149
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_177
timestamp 1644511149
transform 1 0 17388 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1644511149
transform 1 0 19780 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_210
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_216
timestamp 1644511149
transform 1 0 20976 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_232
timestamp 1644511149
transform 1 0 22448 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1644511149
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_252
timestamp 1644511149
transform 1 0 24288 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_258
timestamp 1644511149
transform 1 0 24840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_262
timestamp 1644511149
transform 1 0 25208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 1644511149
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_287
timestamp 1644511149
transform 1 0 27508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_311
timestamp 1644511149
transform 1 0 29716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_321
timestamp 1644511149
transform 1 0 30636 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_327
timestamp 1644511149
transform 1 0 31188 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_357
timestamp 1644511149
transform 1 0 33948 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_362
timestamp 1644511149
transform 1 0 34408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_386
timestamp 1644511149
transform 1 0 36616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_396
timestamp 1644511149
transform 1 0 37536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1644511149
transform 1 0 38180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_101
timestamp 1644511149
transform 1 0 10396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_118
timestamp 1644511149
transform 1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1644511149
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_148
timestamp 1644511149
transform 1 0 14720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1644511149
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1644511149
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1644511149
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_201
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_225
timestamp 1644511149
transform 1 0 21804 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_229
timestamp 1644511149
transform 1 0 22172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_234
timestamp 1644511149
transform 1 0 22632 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_259
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_271
timestamp 1644511149
transform 1 0 26036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_282
timestamp 1644511149
transform 1 0 27048 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_290
timestamp 1644511149
transform 1 0 27784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_323
timestamp 1644511149
transform 1 0 30820 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_331
timestamp 1644511149
transform 1 0 31556 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1644511149
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_350
timestamp 1644511149
transform 1 0 33304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_371
timestamp 1644511149
transform 1 0 35236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_378
timestamp 1644511149
transform 1 0 35880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1644511149
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1644511149
transform 1 0 9200 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1644511149
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_101
timestamp 1644511149
transform 1 0 10396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1644511149
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1644511149
transform 1 0 12420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 1644511149
transform 1 0 13248 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_142
timestamp 1644511149
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1644511149
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_160
timestamp 1644511149
transform 1 0 15824 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_192
timestamp 1644511149
transform 1 0 18768 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_234
timestamp 1644511149
transform 1 0 22632 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_238
timestamp 1644511149
transform 1 0 23000 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1644511149
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1644511149
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_288
timestamp 1644511149
transform 1 0 27600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_302
timestamp 1644511149
transform 1 0 28888 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_330
timestamp 1644511149
transform 1 0 31464 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_348
timestamp 1644511149
transform 1 0 33120 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_357
timestamp 1644511149
transform 1 0 33948 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_365
timestamp 1644511149
transform 1 0 34684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_396
timestamp 1644511149
transform 1 0 37536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1644511149
transform 1 0 38180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_94
timestamp 1644511149
transform 1 0 9752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_98
timestamp 1644511149
transform 1 0 10120 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1644511149
transform 1 0 10856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_120
timestamp 1644511149
transform 1 0 12144 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_164
timestamp 1644511149
transform 1 0 16192 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1644511149
transform 1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_184
timestamp 1644511149
transform 1 0 18032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_220
timestamp 1644511149
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_227
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_241
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_256
timestamp 1644511149
transform 1 0 24656 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_262
timestamp 1644511149
transform 1 0 25208 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_270
timestamp 1644511149
transform 1 0 25944 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_282
timestamp 1644511149
transform 1 0 27048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_290
timestamp 1644511149
transform 1 0 27784 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_317
timestamp 1644511149
transform 1 0 30268 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_329
timestamp 1644511149
transform 1 0 31372 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1644511149
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_344
timestamp 1644511149
transform 1 0 32752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1644511149
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1644511149
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_369
timestamp 1644511149
transform 1 0 35052 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_381
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_9
timestamp 1644511149
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_21
timestamp 1644511149
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_33
timestamp 1644511149
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1644511149
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1644511149
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_91
timestamp 1644511149
transform 1 0 9476 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_99
timestamp 1644511149
transform 1 0 10212 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_120
timestamp 1644511149
transform 1 0 12144 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_133
timestamp 1644511149
transform 1 0 13340 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_139
timestamp 1644511149
transform 1 0 13892 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1644511149
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1644511149
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1644511149
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_176
timestamp 1644511149
transform 1 0 17296 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_210
timestamp 1644511149
transform 1 0 20424 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_216
timestamp 1644511149
transform 1 0 20976 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_245
timestamp 1644511149
transform 1 0 23644 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_253
timestamp 1644511149
transform 1 0 24380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_264
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_285
timestamp 1644511149
transform 1 0 27324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1644511149
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_306
timestamp 1644511149
transform 1 0 29256 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_322
timestamp 1644511149
transform 1 0 30728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1644511149
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_350
timestamp 1644511149
transform 1 0 33304 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_358
timestamp 1644511149
transform 1 0 34040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_380
timestamp 1644511149
transform 1 0 36064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1644511149
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_396
timestamp 1644511149
transform 1 0 37536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_6
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_13
timestamp 1644511149
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1644511149
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_57
timestamp 1644511149
transform 1 0 6348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_61
timestamp 1644511149
transform 1 0 6716 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1644511149
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1644511149
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1644511149
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_95
timestamp 1644511149
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_105
timestamp 1644511149
transform 1 0 10764 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_114
timestamp 1644511149
transform 1 0 11592 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_122
timestamp 1644511149
transform 1 0 12328 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1644511149
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_173
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_186
timestamp 1644511149
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1644511149
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_230
timestamp 1644511149
transform 1 0 22264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1644511149
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1644511149
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_257
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1644511149
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_278
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_287
timestamp 1644511149
transform 1 0 27508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_322
timestamp 1644511149
transform 1 0 30728 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_331
timestamp 1644511149
transform 1 0 31556 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_353
timestamp 1644511149
transform 1 0 33580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1644511149
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_370
timestamp 1644511149
transform 1 0 35144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_73
timestamp 1644511149
transform 1 0 7820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_86
timestamp 1644511149
transform 1 0 9016 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_99
timestamp 1644511149
transform 1 0 10212 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_139
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1644511149
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1644511149
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_185
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1644511149
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1644511149
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_235
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_263
timestamp 1644511149
transform 1 0 25300 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1644511149
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_292
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_299
timestamp 1644511149
transform 1 0 28612 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_310
timestamp 1644511149
transform 1 0 29624 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_324
timestamp 1644511149
transform 1 0 30912 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_344
timestamp 1644511149
transform 1 0 32752 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_353
timestamp 1644511149
transform 1 0 33580 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_364
timestamp 1644511149
transform 1 0 34592 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1644511149
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_397
timestamp 1644511149
transform 1 0 37628 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_57
timestamp 1644511149
transform 1 0 6348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_61
timestamp 1644511149
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1644511149
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_101
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_111
timestamp 1644511149
transform 1 0 11316 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_123
timestamp 1644511149
transform 1 0 12420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_155
timestamp 1644511149
transform 1 0 15364 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_179
timestamp 1644511149
transform 1 0 17572 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1644511149
transform 1 0 18124 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_202
timestamp 1644511149
transform 1 0 19688 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_210
timestamp 1644511149
transform 1 0 20424 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_232
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_238
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_256
timestamp 1644511149
transform 1 0 24656 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1644511149
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_276
timestamp 1644511149
transform 1 0 26496 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1644511149
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_315
timestamp 1644511149
transform 1 0 30084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_335
timestamp 1644511149
transform 1 0 31924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_344
timestamp 1644511149
transform 1 0 32752 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1644511149
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_381
timestamp 1644511149
transform 1 0 36156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1644511149
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 1644511149
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_11
timestamp 1644511149
transform 1 0 2116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_23
timestamp 1644511149
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_35
timestamp 1644511149
transform 1 0 4324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1644511149
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_65
timestamp 1644511149
transform 1 0 7084 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_78
timestamp 1644511149
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_87
timestamp 1644511149
transform 1 0 9108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_95
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1644511149
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1644511149
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_119
timestamp 1644511149
transform 1 0 12052 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_130
timestamp 1644511149
transform 1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_158
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1644511149
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_174
timestamp 1644511149
transform 1 0 17112 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_210
timestamp 1644511149
transform 1 0 20424 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_231
timestamp 1644511149
transform 1 0 22356 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1644511149
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_262
timestamp 1644511149
transform 1 0 25208 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_268
timestamp 1644511149
transform 1 0 25760 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_285
timestamp 1644511149
transform 1 0 27324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1644511149
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_313
timestamp 1644511149
transform 1 0 29900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_324
timestamp 1644511149
transform 1 0 30912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_347
timestamp 1644511149
transform 1 0 33028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_357
timestamp 1644511149
transform 1 0 33948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_364
timestamp 1644511149
transform 1 0 34592 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_397
timestamp 1644511149
transform 1 0 37628 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_8
timestamp 1644511149
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1644511149
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1644511149
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1644511149
transform 1 0 6440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_72
timestamp 1644511149
transform 1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_91
timestamp 1644511149
transform 1 0 9476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1644511149
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp 1644511149
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_119
timestamp 1644511149
transform 1 0 12052 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_128
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_157
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_203
timestamp 1644511149
transform 1 0 19780 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_212
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_238
timestamp 1644511149
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1644511149
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_273
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_300
timestamp 1644511149
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_318
timestamp 1644511149
transform 1 0 30360 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_344
timestamp 1644511149
transform 1 0 32752 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_352
timestamp 1644511149
transform 1 0 33488 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_376
timestamp 1644511149
transform 1 0 35696 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_67
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_79
timestamp 1644511149
transform 1 0 8372 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_103
timestamp 1644511149
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_129
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_140
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_157
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_197
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_235
timestamp 1644511149
transform 1 0 22724 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_246
timestamp 1644511149
transform 1 0 23736 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_252
timestamp 1644511149
transform 1 0 24288 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1644511149
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_260
timestamp 1644511149
transform 1 0 25024 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_265
timestamp 1644511149
transform 1 0 25484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_271
timestamp 1644511149
transform 1 0 26036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_315
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_326
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1644511149
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_340
timestamp 1644511149
transform 1 0 32384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_344
timestamp 1644511149
transform 1 0 32752 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_355
timestamp 1644511149
transform 1 0 33764 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_362
timestamp 1644511149
transform 1 0 34408 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_386
timestamp 1644511149
transform 1 0 36616 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_400
timestamp 1644511149
transform 1 0 37904 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1644511149
transform 1 0 38456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1644511149
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_88
timestamp 1644511149
transform 1 0 9200 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_100
timestamp 1644511149
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_104
timestamp 1644511149
transform 1 0 10672 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_114
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_120
timestamp 1644511149
transform 1 0 12144 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1644511149
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_151
timestamp 1644511149
transform 1 0 14996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1644511149
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_164
timestamp 1644511149
transform 1 0 16192 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1644511149
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_181
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_187
timestamp 1644511149
transform 1 0 18308 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_200
timestamp 1644511149
transform 1 0 19504 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_211
timestamp 1644511149
transform 1 0 20516 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1644511149
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_231
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1644511149
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_261
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_267
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_288
timestamp 1644511149
transform 1 0 27600 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_297
timestamp 1644511149
transform 1 0 28428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_315
timestamp 1644511149
transform 1 0 30084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_339
timestamp 1644511149
transform 1 0 32292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_343
timestamp 1644511149
transform 1 0 32660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_350
timestamp 1644511149
transform 1 0 33304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_354
timestamp 1644511149
transform 1 0 33672 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_373
timestamp 1644511149
transform 1 0 35420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_381
timestamp 1644511149
transform 1 0 36156 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_65
timestamp 1644511149
transform 1 0 7084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_72
timestamp 1644511149
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_76
timestamp 1644511149
transform 1 0 8096 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1644511149
transform 1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_95
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1644511149
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_120
timestamp 1644511149
transform 1 0 12144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_131
timestamp 1644511149
transform 1 0 13156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_141
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_153
timestamp 1644511149
transform 1 0 15180 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_176
timestamp 1644511149
transform 1 0 17296 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1644511149
transform 1 0 17848 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_187
timestamp 1644511149
transform 1 0 18308 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_195
timestamp 1644511149
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_206
timestamp 1644511149
transform 1 0 20056 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_212
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1644511149
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_236
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_244
timestamp 1644511149
transform 1 0 23552 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_266
timestamp 1644511149
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_301
timestamp 1644511149
transform 1 0 28796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_309
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1644511149
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_324
timestamp 1644511149
transform 1 0 30912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_340
timestamp 1644511149
transform 1 0 32384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_347
timestamp 1644511149
transform 1 0 33028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_354
timestamp 1644511149
transform 1 0 33672 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_358
timestamp 1644511149
transform 1 0 34040 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_363
timestamp 1644511149
transform 1 0 34500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_396
timestamp 1644511149
transform 1 0 37536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1644511149
transform 1 0 38180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_61
timestamp 1644511149
transform 1 0 6716 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_79
timestamp 1644511149
transform 1 0 8372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_101
timestamp 1644511149
transform 1 0 10396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_113
timestamp 1644511149
transform 1 0 11500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_124
timestamp 1644511149
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1644511149
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_162
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_170
timestamp 1644511149
transform 1 0 16744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_179
timestamp 1644511149
transform 1 0 17572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_186
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_213
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_234
timestamp 1644511149
transform 1 0 22632 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_242
timestamp 1644511149
transform 1 0 23368 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_260
timestamp 1644511149
transform 1 0 25024 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_267
timestamp 1644511149
transform 1 0 25668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_278
timestamp 1644511149
transform 1 0 26680 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_285
timestamp 1644511149
transform 1 0 27324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_292
timestamp 1644511149
transform 1 0 27968 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_335
timestamp 1644511149
transform 1 0 31924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1644511149
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_375
timestamp 1644511149
transform 1 0 35604 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_402
timestamp 1644511149
transform 1 0 38088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1644511149
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_65
timestamp 1644511149
transform 1 0 7084 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_78
timestamp 1644511149
transform 1 0 8280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1644511149
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_89
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_95
timestamp 1644511149
transform 1 0 9844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_102
timestamp 1644511149
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1644511149
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_121
timestamp 1644511149
transform 1 0 12236 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_143
timestamp 1644511149
transform 1 0 14260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_151
timestamp 1644511149
transform 1 0 14996 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_158
timestamp 1644511149
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1644511149
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_192
timestamp 1644511149
transform 1 0 18768 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_200
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1644511149
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_245
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1644511149
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_267
timestamp 1644511149
transform 1 0 25668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_274
timestamp 1644511149
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_287
timestamp 1644511149
transform 1 0 27508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_299
timestamp 1644511149
transform 1 0 28612 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_311
timestamp 1644511149
transform 1 0 29716 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_319
timestamp 1644511149
transform 1 0 30452 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_326
timestamp 1644511149
transform 1 0 31096 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1644511149
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_346
timestamp 1644511149
transform 1 0 32936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_353
timestamp 1644511149
transform 1 0 33580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_377
timestamp 1644511149
transform 1 0 35788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_381
timestamp 1644511149
transform 1 0 36156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_396
timestamp 1644511149
transform 1 0 37536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1644511149
transform 1 0 38180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_59
timestamp 1644511149
transform 1 0 6532 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_69
timestamp 1644511149
transform 1 0 7452 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1644511149
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_89
timestamp 1644511149
transform 1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_96
timestamp 1644511149
transform 1 0 9936 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_102
timestamp 1644511149
transform 1 0 10488 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_119
timestamp 1644511149
transform 1 0 12052 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1644511149
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_184
timestamp 1644511149
transform 1 0 18032 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_201
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_211
timestamp 1644511149
transform 1 0 20516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_227
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1644511149
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_244
timestamp 1644511149
transform 1 0 23552 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_256
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_262
timestamp 1644511149
transform 1 0 25208 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_268
timestamp 1644511149
transform 1 0 25760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1644511149
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1644511149
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_329
timestamp 1644511149
transform 1 0 31372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_336
timestamp 1644511149
transform 1 0 32016 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_343
timestamp 1644511149
transform 1 0 32660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_350
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_356
timestamp 1644511149
transform 1 0 33856 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_368
timestamp 1644511149
transform 1 0 34960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_375
timestamp 1644511149
transform 1 0 35604 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_381
timestamp 1644511149
transform 1 0 36156 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1644511149
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 1644511149
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_65
timestamp 1644511149
transform 1 0 7084 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_74
timestamp 1644511149
transform 1 0 7912 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_83
timestamp 1644511149
transform 1 0 8740 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_99
timestamp 1644511149
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_121
timestamp 1644511149
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_128
timestamp 1644511149
transform 1 0 12880 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1644511149
transform 1 0 14352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_154
timestamp 1644511149
transform 1 0 15272 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_176
timestamp 1644511149
transform 1 0 17296 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_200
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_208
timestamp 1644511149
transform 1 0 20240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_231
timestamp 1644511149
transform 1 0 22356 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_239
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1644511149
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_284
timestamp 1644511149
transform 1 0 27232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_288
timestamp 1644511149
transform 1 0 27600 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_309
timestamp 1644511149
transform 1 0 29532 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_313
timestamp 1644511149
transform 1 0 29900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_319
timestamp 1644511149
transform 1 0 30452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_357
timestamp 1644511149
transform 1 0 33948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_381
timestamp 1644511149
transform 1 0 36156 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1644511149
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_400
timestamp 1644511149
transform 1 0 37904 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_406
timestamp 1644511149
transform 1 0 38456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1644511149
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_59
timestamp 1644511149
transform 1 0 6532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1644511149
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1644511149
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_108
timestamp 1644511149
transform 1 0 11040 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_124
timestamp 1644511149
transform 1 0 12512 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_157
timestamp 1644511149
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_166
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_174
timestamp 1644511149
transform 1 0 17112 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_179
timestamp 1644511149
transform 1 0 17572 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_183
timestamp 1644511149
transform 1 0 17940 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_187
timestamp 1644511149
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_201
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_227
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_236
timestamp 1644511149
transform 1 0 22816 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1644511149
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_257
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1644511149
transform 1 0 26036 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_281
timestamp 1644511149
transform 1 0 26956 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_290
timestamp 1644511149
transform 1 0 27784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_298
timestamp 1644511149
transform 1 0 28520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1644511149
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_313
timestamp 1644511149
transform 1 0 29900 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_337
timestamp 1644511149
transform 1 0 32108 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_356
timestamp 1644511149
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_368
timestamp 1644511149
transform 1 0 34960 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_375
timestamp 1644511149
transform 1 0 35604 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_381
timestamp 1644511149
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1644511149
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_29
timestamp 1644511149
transform 1 0 3772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_41
timestamp 1644511149
transform 1 0 4876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1644511149
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_65
timestamp 1644511149
transform 1 0 7084 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1644511149
transform 1 0 7544 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_82
timestamp 1644511149
transform 1 0 8648 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_88
timestamp 1644511149
transform 1 0 9200 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_100
timestamp 1644511149
transform 1 0 10304 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_131
timestamp 1644511149
transform 1 0 13156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_139
timestamp 1644511149
transform 1 0 13892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1644511149
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_153
timestamp 1644511149
transform 1 0 15180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_189
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_197
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_203
timestamp 1644511149
transform 1 0 19780 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1644511149
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_234
timestamp 1644511149
transform 1 0 22632 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_238
timestamp 1644511149
transform 1 0 23000 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_245
timestamp 1644511149
transform 1 0 23644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_260
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_267
timestamp 1644511149
transform 1 0 25668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_294
timestamp 1644511149
transform 1 0 28152 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1644511149
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_303
timestamp 1644511149
transform 1 0 28980 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1644511149
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_347
timestamp 1644511149
transform 1 0 33028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_357
timestamp 1644511149
transform 1 0 33948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_381
timestamp 1644511149
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1644511149
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_396
timestamp 1644511149
transform 1 0 37536 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_12
timestamp 1644511149
transform 1 0 2208 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_61
timestamp 1644511149
transform 1 0 6716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_67
timestamp 1644511149
transform 1 0 7268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_90
timestamp 1644511149
transform 1 0 9384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_104
timestamp 1644511149
transform 1 0 10672 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_116
timestamp 1644511149
transform 1 0 11776 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_144
timestamp 1644511149
transform 1 0 14352 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_166
timestamp 1644511149
transform 1 0 16376 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_176
timestamp 1644511149
transform 1 0 17296 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_182
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_218
timestamp 1644511149
transform 1 0 21160 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_225
timestamp 1644511149
transform 1 0 21804 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_229
timestamp 1644511149
transform 1 0 22172 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1644511149
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_258
timestamp 1644511149
transform 1 0 24840 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_266
timestamp 1644511149
transform 1 0 25576 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_278
timestamp 1644511149
transform 1 0 26680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_286
timestamp 1644511149
transform 1 0 27416 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_294
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_323
timestamp 1644511149
transform 1 0 30820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_331
timestamp 1644511149
transform 1 0 31556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_343
timestamp 1644511149
transform 1 0 32660 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_351
timestamp 1644511149
transform 1 0 33396 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_370
timestamp 1644511149
transform 1 0 35144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_393
timestamp 1644511149
transform 1 0 37260 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_400
timestamp 1644511149
transform 1 0 37904 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1644511149
transform 1 0 38456 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_78
timestamp 1644511149
transform 1 0 8280 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1644511149
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_118
timestamp 1644511149
transform 1 0 11960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_130
timestamp 1644511149
transform 1 0 13064 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1644511149
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_174
timestamp 1644511149
transform 1 0 17112 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_185
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_196
timestamp 1644511149
transform 1 0 19136 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_207
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_246
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_270
timestamp 1644511149
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1644511149
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_302
timestamp 1644511149
transform 1 0 28888 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_316
timestamp 1644511149
transform 1 0 30176 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_324
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_342
timestamp 1644511149
transform 1 0 32568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_352
timestamp 1644511149
transform 1 0 33488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_360
timestamp 1644511149
transform 1 0 34224 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_367
timestamp 1644511149
transform 1 0 34868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_374
timestamp 1644511149
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_386
timestamp 1644511149
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_396
timestamp 1644511149
transform 1 0 37536 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_404
timestamp 1644511149
transform 1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_63
timestamp 1644511149
transform 1 0 6900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_74
timestamp 1644511149
transform 1 0 7912 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1644511149
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_96
timestamp 1644511149
transform 1 0 9936 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_104
timestamp 1644511149
transform 1 0 10672 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_144
timestamp 1644511149
transform 1 0 14352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_151
timestamp 1644511149
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_160
timestamp 1644511149
transform 1 0 15824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_170
timestamp 1644511149
transform 1 0 16744 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_178
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1644511149
transform 1 0 18124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_203
timestamp 1644511149
transform 1 0 19780 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_210
timestamp 1644511149
transform 1 0 20424 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_229
timestamp 1644511149
transform 1 0 22172 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_237
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_257
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_268
timestamp 1644511149
transform 1 0 25760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1644511149
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1644511149
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_312
timestamp 1644511149
transform 1 0 29808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_322
timestamp 1644511149
transform 1 0 30728 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_349
timestamp 1644511149
transform 1 0 33212 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_371
timestamp 1644511149
transform 1 0 35236 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_379
timestamp 1644511149
transform 1 0 35972 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1644511149
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_61
timestamp 1644511149
transform 1 0 6716 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_78
timestamp 1644511149
transform 1 0 8280 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_86
timestamp 1644511149
transform 1 0 9016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_94
timestamp 1644511149
transform 1 0 9752 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_101
timestamp 1644511149
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1644511149
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_120
timestamp 1644511149
transform 1 0 12144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_131
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_139
timestamp 1644511149
transform 1 0 13892 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_146
timestamp 1644511149
transform 1 0 14536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_155
timestamp 1644511149
transform 1 0 15364 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1644511149
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_189
timestamp 1644511149
transform 1 0 18492 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_198
timestamp 1644511149
transform 1 0 19320 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_206
timestamp 1644511149
transform 1 0 20056 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_211
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1644511149
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_229
timestamp 1644511149
transform 1 0 22172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_236
timestamp 1644511149
transform 1 0 22816 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_262
timestamp 1644511149
transform 1 0 25208 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_268
timestamp 1644511149
transform 1 0 25760 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_288
timestamp 1644511149
transform 1 0 27600 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_292
timestamp 1644511149
transform 1 0 27968 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_297
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_313
timestamp 1644511149
transform 1 0 29900 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_321
timestamp 1644511149
transform 1 0 30636 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_327
timestamp 1644511149
transform 1 0 31188 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_341
timestamp 1644511149
transform 1 0 32476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_347
timestamp 1644511149
transform 1 0 33028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_359
timestamp 1644511149
transform 1 0 34132 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_383
timestamp 1644511149
transform 1 0 36340 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_400
timestamp 1644511149
transform 1 0 37904 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1644511149
transform 1 0 38456 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_75
timestamp 1644511149
transform 1 0 8004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_90
timestamp 1644511149
transform 1 0 9384 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_98
timestamp 1644511149
transform 1 0 10120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_106
timestamp 1644511149
transform 1 0 10856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_114
timestamp 1644511149
transform 1 0 11592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_120
timestamp 1644511149
transform 1 0 12144 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_128
timestamp 1644511149
transform 1 0 12880 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1644511149
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_161
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_172
timestamp 1644511149
transform 1 0 16928 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_181
timestamp 1644511149
transform 1 0 17756 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1644511149
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_227
timestamp 1644511149
transform 1 0 21988 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_234
timestamp 1644511149
transform 1 0 22632 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_293
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_315
timestamp 1644511149
transform 1 0 30084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_325
timestamp 1644511149
transform 1 0 31004 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_344
timestamp 1644511149
transform 1 0 32752 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_370
timestamp 1644511149
transform 1 0 35144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_381
timestamp 1644511149
transform 1 0 36156 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1644511149
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_64
timestamp 1644511149
transform 1 0 6992 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_73
timestamp 1644511149
transform 1 0 7820 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_79
timestamp 1644511149
transform 1 0 8372 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_83
timestamp 1644511149
transform 1 0 8740 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1644511149
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_121
timestamp 1644511149
transform 1 0 12236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_129
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_135
timestamp 1644511149
transform 1 0 13524 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_139
timestamp 1644511149
transform 1 0 13892 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_150
timestamp 1644511149
transform 1 0 14904 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_156
timestamp 1644511149
transform 1 0 15456 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_177
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_183
timestamp 1644511149
transform 1 0 17940 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_191
timestamp 1644511149
transform 1 0 18676 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_213
timestamp 1644511149
transform 1 0 20700 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_246
timestamp 1644511149
transform 1 0 23736 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_256
timestamp 1644511149
transform 1 0 24656 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_268
timestamp 1644511149
transform 1 0 25760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_288
timestamp 1644511149
transform 1 0 27600 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_294
timestamp 1644511149
transform 1 0 28152 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_312
timestamp 1644511149
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_325
timestamp 1644511149
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_340
timestamp 1644511149
transform 1 0 32384 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_352
timestamp 1644511149
transform 1 0 33488 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_359
timestamp 1644511149
transform 1 0 34132 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_363
timestamp 1644511149
transform 1 0 34500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1644511149
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_399
timestamp 1644511149
transform 1 0 37812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_35
timestamp 1644511149
transform 1 0 4324 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_56
timestamp 1644511149
transform 1 0 6256 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_71
timestamp 1644511149
transform 1 0 7636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_105
timestamp 1644511149
transform 1 0 10764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_117
timestamp 1644511149
transform 1 0 11868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_129
timestamp 1644511149
transform 1 0 12972 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_151
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_159
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_171
timestamp 1644511149
transform 1 0 16836 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_179
timestamp 1644511149
transform 1 0 17572 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_204
timestamp 1644511149
transform 1 0 19872 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_212
timestamp 1644511149
transform 1 0 20608 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_234
timestamp 1644511149
transform 1 0 22632 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_241
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_268
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_276
timestamp 1644511149
transform 1 0 26496 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_282
timestamp 1644511149
transform 1 0 27048 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_293
timestamp 1644511149
transform 1 0 28060 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1644511149
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_323
timestamp 1644511149
transform 1 0 30820 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_336
timestamp 1644511149
transform 1 0 32016 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_352
timestamp 1644511149
transform 1 0 33488 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1644511149
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_370
timestamp 1644511149
transform 1 0 35144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_381
timestamp 1644511149
transform 1 0 36156 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_42
timestamp 1644511149
transform 1 0 4968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_80
timestamp 1644511149
transform 1 0 8464 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_92
timestamp 1644511149
transform 1 0 9568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_102
timestamp 1644511149
transform 1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1644511149
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_117
timestamp 1644511149
transform 1 0 11868 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_128
timestamp 1644511149
transform 1 0 12880 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_141
timestamp 1644511149
transform 1 0 14076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_146
timestamp 1644511149
transform 1 0 14536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1644511149
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_185
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_192
timestamp 1644511149
transform 1 0 18768 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_203
timestamp 1644511149
transform 1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_210
timestamp 1644511149
transform 1 0 20424 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_234
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_241
timestamp 1644511149
transform 1 0 23276 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_250
timestamp 1644511149
transform 1 0 24104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_274
timestamp 1644511149
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_289
timestamp 1644511149
transform 1 0 27692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_296
timestamp 1644511149
transform 1 0 28336 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_307
timestamp 1644511149
transform 1 0 29348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_311
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_341
timestamp 1644511149
transform 1 0 32476 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_356
timestamp 1644511149
transform 1 0 33856 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_380
timestamp 1644511149
transform 1 0 36064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_387
timestamp 1644511149
transform 1 0 36708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_397
timestamp 1644511149
transform 1 0 37628 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_55
timestamp 1644511149
transform 1 0 6164 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_63
timestamp 1644511149
transform 1 0 6900 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_71
timestamp 1644511149
transform 1 0 7636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1644511149
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_96
timestamp 1644511149
transform 1 0 9936 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_102
timestamp 1644511149
transform 1 0 10488 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_118
timestamp 1644511149
transform 1 0 11960 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_124
timestamp 1644511149
transform 1 0 12512 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_172
timestamp 1644511149
transform 1 0 16928 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_180
timestamp 1644511149
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1644511149
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_201
timestamp 1644511149
transform 1 0 19596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_222
timestamp 1644511149
transform 1 0 21528 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1644511149
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_260
timestamp 1644511149
transform 1 0 25024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_284
timestamp 1644511149
transform 1 0 27232 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_292
timestamp 1644511149
transform 1 0 27968 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_300
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_316
timestamp 1644511149
transform 1 0 30176 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_324
timestamp 1644511149
transform 1 0 30912 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_332
timestamp 1644511149
transform 1 0 31648 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1644511149
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_374
timestamp 1644511149
transform 1 0 35512 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1644511149
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_13
timestamp 1644511149
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_25
timestamp 1644511149
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_37
timestamp 1644511149
transform 1 0 4508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_41
timestamp 1644511149
transform 1 0 4876 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_45
timestamp 1644511149
transform 1 0 5244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1644511149
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_63
timestamp 1644511149
transform 1 0 6900 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_76
timestamp 1644511149
transform 1 0 8096 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_86
timestamp 1644511149
transform 1 0 9016 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_95
timestamp 1644511149
transform 1 0 9844 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_104
timestamp 1644511149
transform 1 0 10672 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1644511149
transform 1 0 11960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_142
timestamp 1644511149
transform 1 0 14168 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_150
timestamp 1644511149
transform 1 0 14904 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_159
timestamp 1644511149
transform 1 0 15732 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_176
timestamp 1644511149
transform 1 0 17296 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_186
timestamp 1644511149
transform 1 0 18216 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_198
timestamp 1644511149
transform 1 0 19320 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_214
timestamp 1644511149
transform 1 0 20792 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1644511149
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_245
timestamp 1644511149
transform 1 0 23644 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1644511149
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_264
timestamp 1644511149
transform 1 0 25392 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_286
timestamp 1644511149
transform 1 0 27416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_299
timestamp 1644511149
transform 1 0 28612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_325
timestamp 1644511149
transform 1 0 31004 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_341
timestamp 1644511149
transform 1 0 32476 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_348
timestamp 1644511149
transform 1 0 33120 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_354
timestamp 1644511149
transform 1 0 33672 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_358
timestamp 1644511149
transform 1 0 34040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_365
timestamp 1644511149
transform 1 0 34684 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_374
timestamp 1644511149
transform 1 0 35512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_381
timestamp 1644511149
transform 1 0 36156 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_398
timestamp 1644511149
transform 1 0 37720 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_406
timestamp 1644511149
transform 1 0 38456 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_37
timestamp 1644511149
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_60
timestamp 1644511149
transform 1 0 6624 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_64
timestamp 1644511149
transform 1 0 6992 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_73
timestamp 1644511149
transform 1 0 7820 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1644511149
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_90
timestamp 1644511149
transform 1 0 9384 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_98
timestamp 1644511149
transform 1 0 10120 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_104
timestamp 1644511149
transform 1 0 10672 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_118
timestamp 1644511149
transform 1 0 11960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_125
timestamp 1644511149
transform 1 0 12604 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_135
timestamp 1644511149
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_144
timestamp 1644511149
transform 1 0 14352 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_158
timestamp 1644511149
transform 1 0 15640 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_168
timestamp 1644511149
transform 1 0 16560 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_176
timestamp 1644511149
transform 1 0 17296 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_183
timestamp 1644511149
transform 1 0 17940 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_217
timestamp 1644511149
transform 1 0 21068 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_225
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_229
timestamp 1644511149
transform 1 0 22172 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_242
timestamp 1644511149
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1644511149
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_260
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_268
timestamp 1644511149
transform 1 0 25760 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_276
timestamp 1644511149
transform 1 0 26496 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_284
timestamp 1644511149
transform 1 0 27232 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_290
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_314
timestamp 1644511149
transform 1 0 29992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_337
timestamp 1644511149
transform 1 0 32108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_351
timestamp 1644511149
transform 1 0 33396 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_375
timestamp 1644511149
transform 1 0 35604 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_381
timestamp 1644511149
transform 1 0 36156 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_403
timestamp 1644511149
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_10
timestamp 1644511149
transform 1 0 2024 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_22
timestamp 1644511149
transform 1 0 3128 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_34
timestamp 1644511149
transform 1 0 4232 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_46
timestamp 1644511149
transform 1 0 5336 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_61
timestamp 1644511149
transform 1 0 6716 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_65
timestamp 1644511149
transform 1 0 7084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_89
timestamp 1644511149
transform 1 0 9292 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_101
timestamp 1644511149
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1644511149
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_121
timestamp 1644511149
transform 1 0 12236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_133
timestamp 1644511149
transform 1 0 13340 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_141
timestamp 1644511149
transform 1 0 14076 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_160
timestamp 1644511149
transform 1 0 15824 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_176
timestamp 1644511149
transform 1 0 17296 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_180
timestamp 1644511149
transform 1 0 17664 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_185
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_198
timestamp 1644511149
transform 1 0 19320 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_245
timestamp 1644511149
transform 1 0 23644 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_256
timestamp 1644511149
transform 1 0 24656 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_262
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_267
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1644511149
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_284
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_316
timestamp 1644511149
transform 1 0 30176 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_322
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_330
timestamp 1644511149
transform 1 0 31464 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_346
timestamp 1644511149
transform 1 0 32936 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_350
timestamp 1644511149
transform 1 0 33304 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_371
timestamp 1644511149
transform 1 0 35236 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_377
timestamp 1644511149
transform 1 0 35788 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_381
timestamp 1644511149
transform 1 0 36156 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_388
timestamp 1644511149
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_399
timestamp 1644511149
transform 1 0 37812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_69
timestamp 1644511149
transform 1 0 7452 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_74
timestamp 1644511149
transform 1 0 7912 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1644511149
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_105
timestamp 1644511149
transform 1 0 10764 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_116
timestamp 1644511149
transform 1 0 11776 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_123
timestamp 1644511149
transform 1 0 12420 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_135
timestamp 1644511149
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_144
timestamp 1644511149
transform 1 0 14352 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_152
timestamp 1644511149
transform 1 0 15088 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_176
timestamp 1644511149
transform 1 0 17296 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_184
timestamp 1644511149
transform 1 0 18032 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_204
timestamp 1644511149
transform 1 0 19872 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_215
timestamp 1644511149
transform 1 0 20884 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_228
timestamp 1644511149
transform 1 0 22080 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_237
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_241
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_247
timestamp 1644511149
transform 1 0 23828 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_259
timestamp 1644511149
transform 1 0 24932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_267
timestamp 1644511149
transform 1 0 25668 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_291
timestamp 1644511149
transform 1 0 27876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_317
timestamp 1644511149
transform 1 0 30268 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_329
timestamp 1644511149
transform 1 0 31372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_340
timestamp 1644511149
transform 1 0 32384 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_349
timestamp 1644511149
transform 1 0 33212 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1644511149
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_368
timestamp 1644511149
transform 1 0 34960 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_380
timestamp 1644511149
transform 1 0 36064 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1644511149
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_12
timestamp 1644511149
transform 1 0 2208 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_24
timestamp 1644511149
transform 1 0 3312 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_30
timestamp 1644511149
transform 1 0 3864 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_38
timestamp 1644511149
transform 1 0 4600 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1644511149
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_77
timestamp 1644511149
transform 1 0 8188 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_82
timestamp 1644511149
transform 1 0 8648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_89
timestamp 1644511149
transform 1 0 9292 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_96
timestamp 1644511149
transform 1 0 9936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_106
timestamp 1644511149
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_117
timestamp 1644511149
transform 1 0 11868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_145
timestamp 1644511149
transform 1 0 14444 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 1644511149
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_175
timestamp 1644511149
transform 1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_185
timestamp 1644511149
transform 1 0 18124 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_196
timestamp 1644511149
transform 1 0 19136 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_233
timestamp 1644511149
transform 1 0 22540 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_246
timestamp 1644511149
transform 1 0 23736 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_252
timestamp 1644511149
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_260
timestamp 1644511149
transform 1 0 25024 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1644511149
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_284
timestamp 1644511149
transform 1 0 27232 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_295
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_323
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_340
timestamp 1644511149
transform 1 0 32384 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_351
timestamp 1644511149
transform 1 0 33396 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_363
timestamp 1644511149
transform 1 0 34500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_375
timestamp 1644511149
transform 1 0 35604 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_383
timestamp 1644511149
transform 1 0 36340 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1644511149
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_396
timestamp 1644511149
transform 1 0 37536 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1644511149
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_10
timestamp 1644511149
transform 1 0 2024 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_17
timestamp 1644511149
transform 1 0 2668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_32
timestamp 1644511149
transform 1 0 4048 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_40
timestamp 1644511149
transform 1 0 4784 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_56
timestamp 1644511149
transform 1 0 6256 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_72
timestamp 1644511149
transform 1 0 7728 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_93
timestamp 1644511149
transform 1 0 9660 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_103
timestamp 1644511149
transform 1 0 10580 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_111
timestamp 1644511149
transform 1 0 11316 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_122
timestamp 1644511149
transform 1 0 12328 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_126
timestamp 1644511149
transform 1 0 12696 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_134
timestamp 1644511149
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_146
timestamp 1644511149
transform 1 0 14536 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_154
timestamp 1644511149
transform 1 0 15272 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_175
timestamp 1644511149
transform 1 0 17204 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_183
timestamp 1644511149
transform 1 0 17940 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_217
timestamp 1644511149
transform 1 0 21068 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1644511149
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_267
timestamp 1644511149
transform 1 0 25668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_276
timestamp 1644511149
transform 1 0 26496 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_283
timestamp 1644511149
transform 1 0 27140 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1644511149
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_315
timestamp 1644511149
transform 1 0 30084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_322
timestamp 1644511149
transform 1 0 30728 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_334
timestamp 1644511149
transform 1 0 31832 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_356
timestamp 1644511149
transform 1 0 33856 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_381
timestamp 1644511149
transform 1 0 36156 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_14
timestamp 1644511149
transform 1 0 2392 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_21
timestamp 1644511149
transform 1 0 3036 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_48
timestamp 1644511149
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_77
timestamp 1644511149
transform 1 0 8188 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_100
timestamp 1644511149
transform 1 0 10304 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1644511149
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_121
timestamp 1644511149
transform 1 0 12236 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_130
timestamp 1644511149
transform 1 0 13064 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_146
timestamp 1644511149
transform 1 0 14536 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_159
timestamp 1644511149
transform 1 0 15732 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_177
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_185
timestamp 1644511149
transform 1 0 18124 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_191
timestamp 1644511149
transform 1 0 18676 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_195
timestamp 1644511149
transform 1 0 19044 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_203
timestamp 1644511149
transform 1 0 19780 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_207
timestamp 1644511149
transform 1 0 20148 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_229
timestamp 1644511149
transform 1 0 22172 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_233
timestamp 1644511149
transform 1 0 22540 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_274
timestamp 1644511149
transform 1 0 26312 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_288
timestamp 1644511149
transform 1 0 27600 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_307
timestamp 1644511149
transform 1 0 29348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_311
timestamp 1644511149
transform 1 0 29716 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_340
timestamp 1644511149
transform 1 0 32384 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_348
timestamp 1644511149
transform 1 0 33120 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_363
timestamp 1644511149
transform 1 0 34500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_398
timestamp 1644511149
transform 1 0 37720 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_406
timestamp 1644511149
transform 1 0 38456 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1644511149
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_34
timestamp 1644511149
transform 1 0 4232 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_42
timestamp 1644511149
transform 1 0 4968 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1644511149
transform 1 0 7176 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1644511149
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_105
timestamp 1644511149
transform 1 0 10764 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_116
timestamp 1644511149
transform 1 0 11776 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_120
timestamp 1644511149
transform 1 0 12144 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_129
timestamp 1644511149
transform 1 0 12972 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1644511149
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_144
timestamp 1644511149
transform 1 0 14352 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_159
timestamp 1644511149
transform 1 0 15732 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_169
timestamp 1644511149
transform 1 0 16652 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_181
timestamp 1644511149
transform 1 0 17756 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_190
timestamp 1644511149
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_200
timestamp 1644511149
transform 1 0 19504 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_208
timestamp 1644511149
transform 1 0 20240 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_223
timestamp 1644511149
transform 1 0 21620 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_235
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_243
timestamp 1644511149
transform 1 0 23460 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_257
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_278
timestamp 1644511149
transform 1 0 26680 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_284
timestamp 1644511149
transform 1 0 27232 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_290
timestamp 1644511149
transform 1 0 27784 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_294
timestamp 1644511149
transform 1 0 28152 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_302
timestamp 1644511149
transform 1 0 28888 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_329
timestamp 1644511149
transform 1 0 31372 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_337
timestamp 1644511149
transform 1 0 32108 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_343
timestamp 1644511149
transform 1 0 32660 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_355
timestamp 1644511149
transform 1 0 33764 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_373
timestamp 1644511149
transform 1 0 35420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_378
timestamp 1644511149
transform 1 0 35880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1644511149
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_28
timestamp 1644511149
transform 1 0 3680 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1644511149
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_77
timestamp 1644511149
transform 1 0 8188 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_82
timestamp 1644511149
transform 1 0 8648 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_90
timestamp 1644511149
transform 1 0 9384 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_96
timestamp 1644511149
transform 1 0 9936 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_103
timestamp 1644511149
transform 1 0 10580 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_135
timestamp 1644511149
transform 1 0 13524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_141
timestamp 1644511149
transform 1 0 14076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_150
timestamp 1644511149
transform 1 0 14904 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_157
timestamp 1644511149
transform 1 0 15548 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1644511149
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_204
timestamp 1644511149
transform 1 0 19872 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_228
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_255
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_264
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_286
timestamp 1644511149
transform 1 0 27416 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1644511149
transform 1 0 30360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1644511149
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_340
timestamp 1644511149
transform 1 0 32384 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_347
timestamp 1644511149
transform 1 0 33028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_359
timestamp 1644511149
transform 1 0 34132 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1644511149
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_397
timestamp 1644511149
transform 1 0 37628 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_52
timestamp 1644511149
transform 1 0 5888 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_68
timestamp 1644511149
transform 1 0 7360 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_75
timestamp 1644511149
transform 1 0 8004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_88
timestamp 1644511149
transform 1 0 9200 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_115
timestamp 1644511149
transform 1 0 11684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_119
timestamp 1644511149
transform 1 0 12052 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_123
timestamp 1644511149
transform 1 0 12420 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 1644511149
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_161
timestamp 1644511149
transform 1 0 15916 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_168
timestamp 1644511149
transform 1 0 16560 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_175
timestamp 1644511149
transform 1 0 17204 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_184
timestamp 1644511149
transform 1 0 18032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_188
timestamp 1644511149
transform 1 0 18400 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_218
timestamp 1644511149
transform 1 0 21160 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_234
timestamp 1644511149
transform 1 0 22632 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_241
timestamp 1644511149
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1644511149
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_256
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_263
timestamp 1644511149
transform 1 0 25300 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_267
timestamp 1644511149
transform 1 0 25668 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_300
timestamp 1644511149
transform 1 0 28704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_312
timestamp 1644511149
transform 1 0 29808 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_319
timestamp 1644511149
transform 1 0 30452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_331
timestamp 1644511149
transform 1 0 31556 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_353
timestamp 1644511149
transform 1 0 33580 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_368
timestamp 1644511149
transform 1 0 34960 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_374
timestamp 1644511149
transform 1 0 35512 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_378
timestamp 1644511149
transform 1 0 35880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1644511149
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_26
timestamp 1644511149
transform 1 0 3496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_77
timestamp 1644511149
transform 1 0 8188 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_100
timestamp 1644511149
transform 1 0 10304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_104
timestamp 1644511149
transform 1 0 10672 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_134
timestamp 1644511149
transform 1 0 13432 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_142
timestamp 1644511149
transform 1 0 14168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_175
timestamp 1644511149
transform 1 0 17204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_179
timestamp 1644511149
transform 1 0 17572 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_201
timestamp 1644511149
transform 1 0 19596 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_209
timestamp 1644511149
transform 1 0 20332 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_246
timestamp 1644511149
transform 1 0 23736 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_271
timestamp 1644511149
transform 1 0 26036 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1644511149
transform 1 0 27416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_300
timestamp 1644511149
transform 1 0 28704 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_325
timestamp 1644511149
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1644511149
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1644511149
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_397
timestamp 1644511149
transform 1 0 37628 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_14
timestamp 1644511149
transform 1 0 2392 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1644511149
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_50
timestamp 1644511149
transform 1 0 5704 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_61
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_68
timestamp 1644511149
transform 1 0 7360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_75
timestamp 1644511149
transform 1 0 8004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_90
timestamp 1644511149
transform 1 0 9384 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_104
timestamp 1644511149
transform 1 0 10672 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_134
timestamp 1644511149
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_144
timestamp 1644511149
transform 1 0 14352 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_151
timestamp 1644511149
transform 1 0 14996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_163
timestamp 1644511149
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1644511149
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_176
timestamp 1644511149
transform 1 0 17296 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_183
timestamp 1644511149
transform 1 0 17940 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_220
timestamp 1644511149
transform 1 0 21344 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_228
timestamp 1644511149
transform 1 0 22080 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_246
timestamp 1644511149
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_256
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_332
timestamp 1644511149
transform 1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_340
timestamp 1644511149
transform 1 0 32384 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_348
timestamp 1644511149
transform 1 0 33120 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1644511149
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_388
timestamp 1644511149
transform 1 0 36800 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_396
timestamp 1644511149
transform 1 0 37536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20884 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1260_
timestamp 1644511149
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1261_
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20976 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1263_
timestamp 1644511149
transform -1 0 20976 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19228 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1267_
timestamp 1644511149
transform 1 0 22724 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1268_
timestamp 1644511149
transform -1 0 23644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1269_
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1273_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1274_
timestamp 1644511149
transform 1 0 28060 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1275_
timestamp 1644511149
transform -1 0 28796 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_1  _1276_
timestamp 1644511149
transform -1 0 28336 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1277_
timestamp 1644511149
transform -1 0 23920 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22816 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1279_
timestamp 1644511149
transform -1 0 18768 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1280_
timestamp 1644511149
transform 1 0 16376 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1281_
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1282_
timestamp 1644511149
transform 1 0 14444 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1283_
timestamp 1644511149
transform 1 0 17572 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1284_
timestamp 1644511149
transform 1 0 5336 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1285_
timestamp 1644511149
transform 1 0 9936 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1286_
timestamp 1644511149
transform 1 0 10304 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1287_
timestamp 1644511149
transform -1 0 14536 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1644511149
transform 1 0 10580 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1289_
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1290_
timestamp 1644511149
transform 1 0 20148 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1292_
timestamp 1644511149
transform -1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1294_
timestamp 1644511149
transform 1 0 27048 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1295_
timestamp 1644511149
transform 1 0 26128 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34224 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1297_
timestamp 1644511149
transform -1 0 30360 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1299_
timestamp 1644511149
transform -1 0 35420 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1300_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1301_
timestamp 1644511149
transform 1 0 32752 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1644511149
transform -1 0 35236 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _1303_
timestamp 1644511149
transform -1 0 33764 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1304_
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25668 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1306_
timestamp 1644511149
transform 1 0 29532 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1307_
timestamp 1644511149
transform 1 0 31280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1309_
timestamp 1644511149
transform -1 0 22816 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1310_
timestamp 1644511149
transform -1 0 22356 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1311_
timestamp 1644511149
transform -1 0 18032 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21620 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1313_
timestamp 1644511149
transform -1 0 18768 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1314_
timestamp 1644511149
transform 1 0 13616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1315_
timestamp 1644511149
transform 1 0 10212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1316_
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_1  _1317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10856 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1318_
timestamp 1644511149
transform -1 0 15180 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1319_
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _1320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7084 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1321_
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1322_
timestamp 1644511149
transform 1 0 10764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _1323_
timestamp 1644511149
transform -1 0 16192 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1324_
timestamp 1644511149
transform -1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1326_
timestamp 1644511149
transform -1 0 20056 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1327_
timestamp 1644511149
transform 1 0 24104 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1328_
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_1  _1329_
timestamp 1644511149
transform 1 0 27784 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _1330_
timestamp 1644511149
transform 1 0 31004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1331_
timestamp 1644511149
transform 1 0 25760 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1644511149
transform -1 0 30452 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1333_
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1334_
timestamp 1644511149
transform -1 0 33488 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1335_
timestamp 1644511149
transform -1 0 33488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28612 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1337_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _1338_
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1341_
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1343_
timestamp 1644511149
transform 1 0 16928 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1344_
timestamp 1644511149
transform -1 0 20148 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1345_
timestamp 1644511149
transform -1 0 21068 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1346_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1347_
timestamp 1644511149
transform -1 0 18676 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1348_
timestamp 1644511149
transform 1 0 19412 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1349_
timestamp 1644511149
transform 1 0 18676 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1350_
timestamp 1644511149
transform 1 0 17572 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 1644511149
transform -1 0 21344 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1352_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1353_
timestamp 1644511149
transform 1 0 21068 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1354_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1355_
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1356_
timestamp 1644511149
transform 1 0 23000 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1644511149
transform 1 0 23828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1358_
timestamp 1644511149
transform -1 0 25116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1359_
timestamp 1644511149
transform 1 0 23736 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1360_
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1361_
timestamp 1644511149
transform -1 0 27508 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1362_
timestamp 1644511149
transform -1 0 25024 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1363_
timestamp 1644511149
transform -1 0 16192 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1364_
timestamp 1644511149
transform -1 0 16376 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1365_
timestamp 1644511149
transform 1 0 17940 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1366_
timestamp 1644511149
transform -1 0 18492 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1367_
timestamp 1644511149
transform -1 0 18676 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1368_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1369_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21160 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1371_
timestamp 1644511149
transform -1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1372_
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1373_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1374_
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1375_
timestamp 1644511149
transform -1 0 17940 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1376_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1378_
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1379_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1380_
timestamp 1644511149
transform 1 0 17204 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1381_
timestamp 1644511149
transform -1 0 15272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1383_
timestamp 1644511149
transform 1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1384_
timestamp 1644511149
transform -1 0 18124 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1385_
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1644511149
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1387_
timestamp 1644511149
transform -1 0 20516 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1388_
timestamp 1644511149
transform 1 0 22448 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1389_
timestamp 1644511149
transform 1 0 26128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1390_
timestamp 1644511149
transform 1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1391_
timestamp 1644511149
transform 1 0 17940 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1392_
timestamp 1644511149
transform 1 0 17848 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1393_
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1394_
timestamp 1644511149
transform -1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1395_
timestamp 1644511149
transform 1 0 23552 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1396_
timestamp 1644511149
transform -1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1400_
timestamp 1644511149
transform -1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1401_
timestamp 1644511149
transform 1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1402_
timestamp 1644511149
transform 1 0 20976 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20884 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1405_
timestamp 1644511149
transform -1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _1406_
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1407_
timestamp 1644511149
transform -1 0 24288 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _1408_
timestamp 1644511149
transform -1 0 29992 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1409_
timestamp 1644511149
transform -1 0 23000 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1644511149
transform -1 0 22264 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1411_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23092 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1412_
timestamp 1644511149
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1413_
timestamp 1644511149
transform 1 0 22356 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _1414_
timestamp 1644511149
transform 1 0 22080 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _1415_
timestamp 1644511149
transform -1 0 22448 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1416_
timestamp 1644511149
transform -1 0 19596 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19688 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18768 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1419_
timestamp 1644511149
transform 1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1420_
timestamp 1644511149
transform 1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1421_
timestamp 1644511149
transform 1 0 16836 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1422_
timestamp 1644511149
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1644511149
transform -1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1424_
timestamp 1644511149
transform 1 0 17020 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1425_
timestamp 1644511149
transform -1 0 19044 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1426_
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1427_
timestamp 1644511149
transform -1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1428_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1429_
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1430_
timestamp 1644511149
transform -1 0 15640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1431_
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1432_
timestamp 1644511149
transform -1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1433_
timestamp 1644511149
transform -1 0 22816 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1434_
timestamp 1644511149
transform -1 0 21252 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _1435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1436_
timestamp 1644511149
transform 1 0 19044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1438_
timestamp 1644511149
transform -1 0 19872 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1439_
timestamp 1644511149
transform 1 0 16836 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1440_
timestamp 1644511149
transform 1 0 17664 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1441_
timestamp 1644511149
transform 1 0 17296 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1442_
timestamp 1644511149
transform -1 0 16468 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1443_
timestamp 1644511149
transform -1 0 19596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1444_
timestamp 1644511149
transform -1 0 19872 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 1644511149
transform 1 0 15364 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1644511149
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1447_
timestamp 1644511149
transform 1 0 16744 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1449_
timestamp 1644511149
transform 1 0 18216 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1451_
timestamp 1644511149
transform 1 0 24656 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1452_
timestamp 1644511149
transform -1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1453_
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1454_
timestamp 1644511149
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1455_
timestamp 1644511149
transform 1 0 25944 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1456_
timestamp 1644511149
transform -1 0 25392 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1457_
timestamp 1644511149
transform -1 0 24196 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1458_
timestamp 1644511149
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1459_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1460_
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1644511149
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1462_
timestamp 1644511149
transform 1 0 22816 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1463_
timestamp 1644511149
transform -1 0 26496 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a31oi_1  _1464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25208 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1465_
timestamp 1644511149
transform -1 0 25760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1467_
timestamp 1644511149
transform -1 0 26404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1468_
timestamp 1644511149
transform 1 0 23460 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1469_
timestamp 1644511149
transform 1 0 24932 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1470_
timestamp 1644511149
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1471_
timestamp 1644511149
transform 1 0 27876 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1472_
timestamp 1644511149
transform 1 0 27968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1473_
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1474_
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1476_
timestamp 1644511149
transform -1 0 27048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1477_
timestamp 1644511149
transform 1 0 27416 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1478_
timestamp 1644511149
transform -1 0 26496 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1479_
timestamp 1644511149
transform -1 0 27600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1480_
timestamp 1644511149
transform -1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1481_
timestamp 1644511149
transform -1 0 26496 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1482_
timestamp 1644511149
transform -1 0 27968 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1483_
timestamp 1644511149
transform 1 0 30176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1484_
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1485_
timestamp 1644511149
transform -1 0 30084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1486_
timestamp 1644511149
transform -1 0 26496 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1487_
timestamp 1644511149
transform 1 0 24104 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1488_
timestamp 1644511149
transform 1 0 25668 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1489_
timestamp 1644511149
transform -1 0 25484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1490_
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1491_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1492_
timestamp 1644511149
transform 1 0 21528 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1493_
timestamp 1644511149
transform 1 0 25392 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1494_
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1496_
timestamp 1644511149
transform -1 0 24288 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1497_
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1498_
timestamp 1644511149
transform -1 0 26220 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1499_
timestamp 1644511149
transform 1 0 27692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1500_
timestamp 1644511149
transform -1 0 26128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1501_
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1502_
timestamp 1644511149
transform -1 0 25576 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1503_
timestamp 1644511149
transform -1 0 25116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1504_
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 1644511149
transform 1 0 20424 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22816 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1507_
timestamp 1644511149
transform -1 0 23644 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1508_
timestamp 1644511149
transform 1 0 23184 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1644511149
transform -1 0 21804 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1510_
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1511_
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1644511149
transform 1 0 20148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1513_
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1514_
timestamp 1644511149
transform 1 0 20424 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _1515_
timestamp 1644511149
transform -1 0 23460 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1516_
timestamp 1644511149
transform -1 0 22632 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1517_
timestamp 1644511149
transform 1 0 16744 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1518_
timestamp 1644511149
transform -1 0 21344 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1519_
timestamp 1644511149
transform 1 0 20792 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _1520_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1521_
timestamp 1644511149
transform 1 0 22264 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1522_
timestamp 1644511149
transform -1 0 23368 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1523_
timestamp 1644511149
transform 1 0 27968 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1524_
timestamp 1644511149
transform 1 0 28888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1525_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1526_
timestamp 1644511149
transform 1 0 30176 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1527_
timestamp 1644511149
transform -1 0 35144 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1528_
timestamp 1644511149
transform -1 0 34684 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1529_
timestamp 1644511149
transform -1 0 33856 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1530_
timestamp 1644511149
transform 1 0 31096 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1644511149
transform -1 0 27968 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1532_
timestamp 1644511149
transform -1 0 29164 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1533_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1534_
timestamp 1644511149
transform 1 0 30452 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1535_
timestamp 1644511149
transform -1 0 35696 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1536_
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1537_
timestamp 1644511149
transform 1 0 32660 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1538_
timestamp 1644511149
transform 1 0 33120 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1539_
timestamp 1644511149
transform -1 0 32568 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1540_
timestamp 1644511149
transform -1 0 31648 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1541_
timestamp 1644511149
transform 1 0 25300 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1542_
timestamp 1644511149
transform 1 0 25208 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1543_
timestamp 1644511149
transform -1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1544_
timestamp 1644511149
transform -1 0 26312 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1545_
timestamp 1644511149
transform -1 0 26220 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1546_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1547_
timestamp 1644511149
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1548_
timestamp 1644511149
transform -1 0 27324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1549_
timestamp 1644511149
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1551_
timestamp 1644511149
transform -1 0 25392 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1552_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1553_
timestamp 1644511149
transform -1 0 26496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1554_
timestamp 1644511149
transform -1 0 26036 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1556_
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1557_
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1558_
timestamp 1644511149
transform -1 0 25944 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1559_
timestamp 1644511149
transform -1 0 32936 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1560_
timestamp 1644511149
transform -1 0 31648 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1561_
timestamp 1644511149
transform -1 0 33120 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1562_
timestamp 1644511149
transform -1 0 32752 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1563_
timestamp 1644511149
transform -1 0 33580 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1564_
timestamp 1644511149
transform -1 0 32384 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _1565_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1566_
timestamp 1644511149
transform 1 0 32108 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1567_
timestamp 1644511149
transform -1 0 31280 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1568_
timestamp 1644511149
transform 1 0 25576 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1569_
timestamp 1644511149
transform 1 0 35052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1570_
timestamp 1644511149
transform 1 0 28980 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1571_
timestamp 1644511149
transform -1 0 30820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30084 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1573_
timestamp 1644511149
transform 1 0 27140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1574_
timestamp 1644511149
transform 1 0 26680 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1575_
timestamp 1644511149
transform 1 0 28152 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1576_
timestamp 1644511149
transform -1 0 28520 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1577_
timestamp 1644511149
transform 1 0 27416 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1578_
timestamp 1644511149
transform -1 0 28152 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1580_
timestamp 1644511149
transform -1 0 31372 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1581_
timestamp 1644511149
transform -1 0 30084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1582_
timestamp 1644511149
transform -1 0 29808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1583_
timestamp 1644511149
transform -1 0 31372 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1584_
timestamp 1644511149
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29992 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1586_
timestamp 1644511149
transform -1 0 31556 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1644511149
transform -1 0 32568 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1588_
timestamp 1644511149
transform -1 0 31648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1589_
timestamp 1644511149
transform -1 0 32568 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1590_
timestamp 1644511149
transform -1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1592_
timestamp 1644511149
transform -1 0 31740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1593_
timestamp 1644511149
transform -1 0 34040 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1594_
timestamp 1644511149
transform 1 0 33304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1595_
timestamp 1644511149
transform 1 0 32476 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1596_
timestamp 1644511149
transform -1 0 35880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1597_
timestamp 1644511149
transform -1 0 35420 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1598_
timestamp 1644511149
transform -1 0 35788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34408 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1600_
timestamp 1644511149
transform -1 0 36064 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1601_
timestamp 1644511149
transform -1 0 35604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1602_
timestamp 1644511149
transform -1 0 34408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1603_
timestamp 1644511149
transform 1 0 35604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1604_
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1605_
timestamp 1644511149
transform 1 0 32660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1606_
timestamp 1644511149
transform 1 0 32292 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1607_
timestamp 1644511149
transform -1 0 33304 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1608_
timestamp 1644511149
transform 1 0 33672 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1609_
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1610_
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1611_
timestamp 1644511149
transform 1 0 33212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1612_
timestamp 1644511149
transform 1 0 29900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1613_
timestamp 1644511149
transform -1 0 33672 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1614_
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1615_
timestamp 1644511149
transform -1 0 32844 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1616_
timestamp 1644511149
transform 1 0 33488 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1617_
timestamp 1644511149
transform -1 0 37536 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1618_
timestamp 1644511149
transform -1 0 34592 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1619_
timestamp 1644511149
transform -1 0 34224 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1620_
timestamp 1644511149
transform 1 0 31280 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1621_
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1622_
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1623_
timestamp 1644511149
transform -1 0 34500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1624_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1625_
timestamp 1644511149
transform -1 0 34592 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1627_
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1628_
timestamp 1644511149
transform -1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1629_
timestamp 1644511149
transform -1 0 30912 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1630_
timestamp 1644511149
transform -1 0 31556 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1631_
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1632_
timestamp 1644511149
transform 1 0 29992 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1633_
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1634_
timestamp 1644511149
transform -1 0 32384 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1635_
timestamp 1644511149
transform -1 0 32752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1636_
timestamp 1644511149
transform -1 0 31372 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1637_
timestamp 1644511149
transform 1 0 33396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1638_
timestamp 1644511149
transform -1 0 27508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1639_
timestamp 1644511149
transform -1 0 31556 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1640_
timestamp 1644511149
transform -1 0 29624 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1641_
timestamp 1644511149
transform -1 0 30728 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1642_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1643_
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1644_
timestamp 1644511149
transform -1 0 29532 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1645_
timestamp 1644511149
transform -1 0 29072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1646_
timestamp 1644511149
transform -1 0 28428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1647_
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1648_
timestamp 1644511149
transform 1 0 28336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1649_
timestamp 1644511149
transform 1 0 27416 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1650_
timestamp 1644511149
transform -1 0 27692 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1644511149
transform -1 0 27324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1652_
timestamp 1644511149
transform 1 0 25576 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1653_
timestamp 1644511149
transform -1 0 26496 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1654_
timestamp 1644511149
transform -1 0 27416 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1655_
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1656_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1657_
timestamp 1644511149
transform -1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1658_
timestamp 1644511149
transform -1 0 23276 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1659_
timestamp 1644511149
transform -1 0 24656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1660_
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1661_
timestamp 1644511149
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1662_
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1663_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1664_
timestamp 1644511149
transform 1 0 18400 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1665_
timestamp 1644511149
transform -1 0 25024 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1666_
timestamp 1644511149
transform -1 0 23920 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1667_
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1668_
timestamp 1644511149
transform 1 0 17020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1669_
timestamp 1644511149
transform 1 0 21160 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand4b_1  _1670_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22080 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _1671_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1672_
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22540 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_4  _1674_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23828 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1675_
timestamp 1644511149
transform -1 0 15640 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1676_
timestamp 1644511149
transform 1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1677_
timestamp 1644511149
transform 1 0 20792 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1678_
timestamp 1644511149
transform -1 0 19044 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1679_
timestamp 1644511149
transform -1 0 11960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1680_
timestamp 1644511149
transform -1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1681_
timestamp 1644511149
transform 1 0 15088 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1682_
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1683_
timestamp 1644511149
transform -1 0 14536 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1684_
timestamp 1644511149
transform 1 0 11040 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1685_
timestamp 1644511149
transform 1 0 6532 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1644511149
transform -1 0 6900 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1687_
timestamp 1644511149
transform 1 0 6992 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1688_
timestamp 1644511149
transform -1 0 11040 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1689_
timestamp 1644511149
transform -1 0 9936 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1690_
timestamp 1644511149
transform 1 0 9384 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1691_
timestamp 1644511149
transform 1 0 11500 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1693_
timestamp 1644511149
transform 1 0 12328 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1694_
timestamp 1644511149
transform 1 0 15548 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1695_
timestamp 1644511149
transform -1 0 18676 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1696_
timestamp 1644511149
transform 1 0 16744 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1697_
timestamp 1644511149
transform -1 0 18768 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1698_
timestamp 1644511149
transform -1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1699_
timestamp 1644511149
transform -1 0 10120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1700_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1701_
timestamp 1644511149
transform 1 0 18492 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1702_
timestamp 1644511149
transform -1 0 18768 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1703_
timestamp 1644511149
transform -1 0 15088 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1704_
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1705_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1706_
timestamp 1644511149
transform 1 0 17296 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1707_
timestamp 1644511149
transform 1 0 17664 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1708_
timestamp 1644511149
transform 1 0 17664 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1709_
timestamp 1644511149
transform -1 0 19320 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1710_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1711_
timestamp 1644511149
transform -1 0 22816 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1712_
timestamp 1644511149
transform -1 0 21344 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1713_
timestamp 1644511149
transform -1 0 17296 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1714_
timestamp 1644511149
transform -1 0 17388 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1715_
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1716_
timestamp 1644511149
transform 1 0 18032 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1717_
timestamp 1644511149
transform 1 0 19136 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1718_
timestamp 1644511149
transform 1 0 19044 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1719_
timestamp 1644511149
transform 1 0 13248 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _1720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17388 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1721_
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1722_
timestamp 1644511149
transform -1 0 19136 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1723_
timestamp 1644511149
transform -1 0 20424 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1724_
timestamp 1644511149
transform -1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1725_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1726_
timestamp 1644511149
transform -1 0 19320 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1728_
timestamp 1644511149
transform -1 0 18308 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1729_
timestamp 1644511149
transform 1 0 19504 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1730_
timestamp 1644511149
transform 1 0 17664 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1731_
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1733_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1734_
timestamp 1644511149
transform -1 0 17296 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1735_
timestamp 1644511149
transform 1 0 15916 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1736_
timestamp 1644511149
transform -1 0 16744 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1737_
timestamp 1644511149
transform -1 0 17756 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1738_
timestamp 1644511149
transform -1 0 16928 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1739_
timestamp 1644511149
transform 1 0 16652 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1740_
timestamp 1644511149
transform -1 0 15364 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1741_
timestamp 1644511149
transform 1 0 15364 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1742_
timestamp 1644511149
transform -1 0 17112 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1743_
timestamp 1644511149
transform -1 0 21344 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1744_
timestamp 1644511149
transform -1 0 15916 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 1644511149
transform 1 0 15548 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1746_
timestamp 1644511149
transform -1 0 14352 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1747_
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1748_
timestamp 1644511149
transform -1 0 15180 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1750_
timestamp 1644511149
transform -1 0 14536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1751_
timestamp 1644511149
transform -1 0 13892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1752_
timestamp 1644511149
transform 1 0 14260 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1753_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp 1644511149
transform -1 0 15732 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1755_
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1756_
timestamp 1644511149
transform 1 0 14904 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1644511149
transform -1 0 14352 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1758_
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1759_
timestamp 1644511149
transform -1 0 12880 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1760_
timestamp 1644511149
transform 1 0 12604 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1761_
timestamp 1644511149
transform -1 0 13340 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1762_
timestamp 1644511149
transform 1 0 12972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1763_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1764_
timestamp 1644511149
transform 1 0 12512 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1765_
timestamp 1644511149
transform -1 0 12144 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1766_
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1767_
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1768_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1769_
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1770_
timestamp 1644511149
transform -1 0 8464 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1771_
timestamp 1644511149
transform -1 0 10672 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1772_
timestamp 1644511149
transform -1 0 8464 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1773_
timestamp 1644511149
transform 1 0 7360 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1774_
timestamp 1644511149
transform -1 0 9384 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1775_
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1776_
timestamp 1644511149
transform 1 0 9292 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1777_
timestamp 1644511149
transform 1 0 9752 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1644511149
transform 1 0 7636 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1779_
timestamp 1644511149
transform 1 0 6992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1780_
timestamp 1644511149
transform 1 0 9108 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1781_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1782_
timestamp 1644511149
transform 1 0 10396 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1783_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1784_
timestamp 1644511149
transform -1 0 7912 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1785_
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1786_
timestamp 1644511149
transform -1 0 7636 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1787_
timestamp 1644511149
transform -1 0 9384 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1788_
timestamp 1644511149
transform -1 0 5888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1789_
timestamp 1644511149
transform 1 0 6808 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1790_
timestamp 1644511149
transform -1 0 8464 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1791_
timestamp 1644511149
transform -1 0 7912 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1792_
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1793_
timestamp 1644511149
transform 1 0 12144 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1794_
timestamp 1644511149
transform -1 0 12604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1795_
timestamp 1644511149
transform -1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1797_
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1798_
timestamp 1644511149
transform 1 0 10212 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1799_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1800_
timestamp 1644511149
transform -1 0 9936 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1801_
timestamp 1644511149
transform -1 0 14352 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1802_
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1803_
timestamp 1644511149
transform 1 0 15272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1804_
timestamp 1644511149
transform -1 0 11776 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1805_
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1806_
timestamp 1644511149
transform 1 0 10672 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1807_
timestamp 1644511149
transform -1 0 12328 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1808_
timestamp 1644511149
transform 1 0 12788 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1809_
timestamp 1644511149
transform 1 0 12788 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1810_
timestamp 1644511149
transform -1 0 13248 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1811_
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1813_
timestamp 1644511149
transform 1 0 15088 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1814_
timestamp 1644511149
transform -1 0 14904 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1815_
timestamp 1644511149
transform -1 0 17296 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1816_
timestamp 1644511149
transform -1 0 15824 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1817_
timestamp 1644511149
transform 1 0 18124 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1818_
timestamp 1644511149
transform -1 0 17756 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 1644511149
transform -1 0 15824 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1820_
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1821_
timestamp 1644511149
transform -1 0 28980 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1822_
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1823_
timestamp 1644511149
transform 1 0 22080 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1824_
timestamp 1644511149
transform 1 0 28796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1825_
timestamp 1644511149
transform -1 0 25760 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1826_
timestamp 1644511149
transform -1 0 23920 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1827_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _1828_
timestamp 1644511149
transform 1 0 31004 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1829_
timestamp 1644511149
transform -1 0 35144 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1830_
timestamp 1644511149
transform -1 0 35144 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1831_
timestamp 1644511149
transform -1 0 32844 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1832_
timestamp 1644511149
transform -1 0 32752 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1833_
timestamp 1644511149
transform -1 0 32384 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1834_
timestamp 1644511149
transform 1 0 30820 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1835_
timestamp 1644511149
transform -1 0 28888 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1836_
timestamp 1644511149
transform -1 0 28704 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1837_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1838_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1839_
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1840_
timestamp 1644511149
transform -1 0 28152 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1841_
timestamp 1644511149
transform 1 0 26772 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1842_
timestamp 1644511149
transform 1 0 26128 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1843_
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1844_
timestamp 1644511149
transform -1 0 31556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1845_
timestamp 1644511149
transform -1 0 26496 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1846_
timestamp 1644511149
transform 1 0 27140 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1847_
timestamp 1644511149
transform -1 0 27784 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1848_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1849_
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1850_
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1851_
timestamp 1644511149
transform 1 0 25484 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1852_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1853_
timestamp 1644511149
transform 1 0 26404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1854_
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1855_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1856_
timestamp 1644511149
transform 1 0 24748 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1857_
timestamp 1644511149
transform 1 0 32292 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1858_
timestamp 1644511149
transform -1 0 33028 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1859_
timestamp 1644511149
transform -1 0 29072 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1860_
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1861_
timestamp 1644511149
transform -1 0 29348 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1862_
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1863_
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1864_
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1865_
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 1644511149
transform -1 0 28060 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1867_
timestamp 1644511149
transform -1 0 27600 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1868_
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1869_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1870_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1871_
timestamp 1644511149
transform 1 0 27324 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1872_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1873_
timestamp 1644511149
transform 1 0 27416 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1874_
timestamp 1644511149
transform -1 0 28888 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1875_
timestamp 1644511149
transform -1 0 24932 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1876_
timestamp 1644511149
transform -1 0 24656 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1877_
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1878_
timestamp 1644511149
transform -1 0 22172 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1879_
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1880_
timestamp 1644511149
transform 1 0 22356 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1881_
timestamp 1644511149
transform -1 0 23828 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1882_
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1883_
timestamp 1644511149
transform -1 0 21344 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1884_
timestamp 1644511149
transform -1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1885_
timestamp 1644511149
transform -1 0 24840 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1886_
timestamp 1644511149
transform 1 0 25300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1887_
timestamp 1644511149
transform -1 0 22540 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1888_
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1889_
timestamp 1644511149
transform 1 0 22264 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1890_
timestamp 1644511149
transform -1 0 25024 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1891_
timestamp 1644511149
transform -1 0 25668 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1892_
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1893_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1894_
timestamp 1644511149
transform -1 0 32660 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1895_
timestamp 1644511149
transform -1 0 32476 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1896_
timestamp 1644511149
transform -1 0 30176 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1897_
timestamp 1644511149
transform 1 0 28612 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1898_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1899_
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1900_
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1901_
timestamp 1644511149
transform 1 0 33764 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1902_
timestamp 1644511149
transform 1 0 33764 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1903_
timestamp 1644511149
transform 1 0 32200 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1904_
timestamp 1644511149
transform -1 0 34224 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1905_
timestamp 1644511149
transform -1 0 33120 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1906_
timestamp 1644511149
transform 1 0 32752 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1907_
timestamp 1644511149
transform 1 0 32200 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1908_
timestamp 1644511149
transform -1 0 28060 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1909_
timestamp 1644511149
transform 1 0 27140 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1910_
timestamp 1644511149
transform -1 0 29348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1911_
timestamp 1644511149
transform 1 0 28428 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1912_
timestamp 1644511149
transform 1 0 28244 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1913_
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1914_
timestamp 1644511149
transform -1 0 27784 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1915_
timestamp 1644511149
transform 1 0 27140 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1916_
timestamp 1644511149
transform 1 0 25392 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1917_
timestamp 1644511149
transform -1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1918_
timestamp 1644511149
transform 1 0 25484 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1919_
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1920_
timestamp 1644511149
transform 1 0 27600 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1921_
timestamp 1644511149
transform 1 0 26036 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1922_
timestamp 1644511149
transform 1 0 26864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1923_
timestamp 1644511149
transform -1 0 32384 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1924_
timestamp 1644511149
transform 1 0 30452 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1925_
timestamp 1644511149
transform -1 0 31648 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1926_
timestamp 1644511149
transform -1 0 30176 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1927_
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1928_
timestamp 1644511149
transform 1 0 33212 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1929_
timestamp 1644511149
transform 1 0 30084 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1930_
timestamp 1644511149
transform -1 0 30084 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1931_
timestamp 1644511149
transform -1 0 32016 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1932_
timestamp 1644511149
transform 1 0 33856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1933_
timestamp 1644511149
transform 1 0 33856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1934_
timestamp 1644511149
transform 1 0 35512 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1935_
timestamp 1644511149
transform -1 0 33856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1936_
timestamp 1644511149
transform 1 0 33764 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1937_
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1938_
timestamp 1644511149
transform -1 0 34224 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1939_
timestamp 1644511149
transform 1 0 34592 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1940_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1941_
timestamp 1644511149
transform -1 0 34132 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1942_
timestamp 1644511149
transform 1 0 35512 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1943_
timestamp 1644511149
transform 1 0 33396 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1944_
timestamp 1644511149
transform 1 0 35236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1945_
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1946_
timestamp 1644511149
transform -1 0 32936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1947_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1948_
timestamp 1644511149
transform -1 0 33856 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1949_
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1950_
timestamp 1644511149
transform -1 0 30268 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1951_
timestamp 1644511149
transform -1 0 31740 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1952_
timestamp 1644511149
transform 1 0 31924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1953_
timestamp 1644511149
transform -1 0 31188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1954_
timestamp 1644511149
transform -1 0 30728 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1955_
timestamp 1644511149
transform -1 0 30820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1956_
timestamp 1644511149
transform 1 0 29624 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1957_
timestamp 1644511149
transform 1 0 29440 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1958_
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1959_
timestamp 1644511149
transform 1 0 28336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1960_
timestamp 1644511149
transform -1 0 6716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _1961_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _1962_
timestamp 1644511149
transform 1 0 33396 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1963_
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1964_
timestamp 1644511149
transform -1 0 2392 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1965_
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1966_
timestamp 1644511149
transform -1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1967_
timestamp 1644511149
transform 1 0 34776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1968_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1969_
timestamp 1644511149
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1970_
timestamp 1644511149
transform 1 0 37904 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1971_
timestamp 1644511149
transform -1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1972_
timestamp 1644511149
transform -1 0 37628 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1973_
timestamp 1644511149
transform -1 0 37536 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1974_
timestamp 1644511149
transform 1 0 4416 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _1975_
timestamp 1644511149
transform 1 0 5152 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1976_
timestamp 1644511149
transform 1 0 37444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1977_
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1978_
timestamp 1644511149
transform 1 0 37352 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1979_
timestamp 1644511149
transform -1 0 4692 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1980_
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1981_
timestamp 1644511149
transform -1 0 5980 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 1644511149
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1983_
timestamp 1644511149
transform 1 0 37536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 1644511149
transform 1 0 37536 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1985_
timestamp 1644511149
transform 1 0 3956 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1986_
timestamp 1644511149
transform 1 0 37628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1987_
timestamp 1644511149
transform 1 0 6624 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1988_
timestamp 1644511149
transform -1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1989_
timestamp 1644511149
transform 1 0 37444 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1990_
timestamp 1644511149
transform -1 0 24656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1991_
timestamp 1644511149
transform -1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1992_
timestamp 1644511149
transform 1 0 37444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1993_
timestamp 1644511149
transform -1 0 5980 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1994_
timestamp 1644511149
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1995_
timestamp 1644511149
transform 1 0 35052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1996_
timestamp 1644511149
transform -1 0 3036 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1997_
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1998_
timestamp 1644511149
transform -1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1999_
timestamp 1644511149
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2000_
timestamp 1644511149
transform 1 0 37352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2001_
timestamp 1644511149
transform 1 0 37352 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2002_
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2003_
timestamp 1644511149
transform -1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2004_
timestamp 1644511149
transform -1 0 4048 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2005_
timestamp 1644511149
transform 1 0 19412 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _2006_
timestamp 1644511149
transform -1 0 21988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2007_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2008_
timestamp 1644511149
transform 1 0 17756 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2009_
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2010_
timestamp 1644511149
transform -1 0 2852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2011_
timestamp 1644511149
transform -1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _2012_
timestamp 1644511149
transform 1 0 22356 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2013_
timestamp 1644511149
transform -1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2014_
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2015_
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2016_
timestamp 1644511149
transform -1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2017_
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2018_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2019_
timestamp 1644511149
transform -1 0 37536 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2020_
timestamp 1644511149
transform -1 0 22172 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2021_
timestamp 1644511149
transform 1 0 37904 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2022_
timestamp 1644511149
transform 1 0 36248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2023_
timestamp 1644511149
transform -1 0 36800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _2024_
timestamp 1644511149
transform 1 0 20884 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2025_
timestamp 1644511149
transform -1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2026_
timestamp 1644511149
transform -1 0 32384 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2027_
timestamp 1644511149
transform -1 0 2300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2028_
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2029_
timestamp 1644511149
transform 1 0 37904 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _2030_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _2031_
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2032_
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2033_
timestamp 1644511149
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2034_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2035_
timestamp 1644511149
transform -1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2036_
timestamp 1644511149
transform 1 0 19504 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _2037_
timestamp 1644511149
transform 1 0 20240 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2038_
timestamp 1644511149
transform 1 0 37444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2039_
timestamp 1644511149
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2040_
timestamp 1644511149
transform -1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2041_
timestamp 1644511149
transform -1 0 2392 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2042_
timestamp 1644511149
transform -1 0 36800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _2043_
timestamp 1644511149
transform -1 0 21344 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2044_
timestamp 1644511149
transform -1 0 37812 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2045_
timestamp 1644511149
transform -1 0 37720 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2046_
timestamp 1644511149
transform -1 0 17204 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2047_
timestamp 1644511149
transform 1 0 37904 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2048_
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _2049_
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2050_
timestamp 1644511149
transform -1 0 33028 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2051_
timestamp 1644511149
transform -1 0 19780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2052_
timestamp 1644511149
transform 1 0 37352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2053_
timestamp 1644511149
transform -1 0 2944 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2054_
timestamp 1644511149
transform 1 0 37444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _2055_
timestamp 1644511149
transform -1 0 21344 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2056_
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2057_
timestamp 1644511149
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2058_
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2059_
timestamp 1644511149
transform -1 0 2668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2060_
timestamp 1644511149
transform 1 0 37904 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _2061_
timestamp 1644511149
transform 1 0 21528 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2062_
timestamp 1644511149
transform -1 0 37812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2063_
timestamp 1644511149
transform -1 0 36800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2064_
timestamp 1644511149
transform -1 0 10672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2065_
timestamp 1644511149
transform -1 0 10580 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2066_
timestamp 1644511149
transform 1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _2067_
timestamp 1644511149
transform 1 0 6256 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2068_
timestamp 1644511149
transform 1 0 10488 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2069_
timestamp 1644511149
transform 1 0 27784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2070_
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2071_
timestamp 1644511149
transform 1 0 37904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2072_
timestamp 1644511149
transform -1 0 3036 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _2073_
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2074_
timestamp 1644511149
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2075_
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2076_
timestamp 1644511149
transform -1 0 22080 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2077_
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2078_
timestamp 1644511149
transform -1 0 36800 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _2079_
timestamp 1644511149
transform -1 0 5888 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2080_
timestamp 1644511149
transform -1 0 23092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2081_
timestamp 1644511149
transform -1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2082_
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2083_
timestamp 1644511149
transform -1 0 7360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2084_
timestamp 1644511149
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _2085_
timestamp 1644511149
transform 1 0 6348 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2086_
timestamp 1644511149
transform -1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2087_
timestamp 1644511149
transform 1 0 34960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2088_
timestamp 1644511149
transform -1 0 9200 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2089_
timestamp 1644511149
transform -1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2090_
timestamp 1644511149
transform -1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2091_
timestamp 1644511149
transform -1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2092_
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2093_
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2094_
timestamp 1644511149
transform -1 0 20884 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2095_
timestamp 1644511149
transform -1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2096_
timestamp 1644511149
transform -1 0 11592 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2097_
timestamp 1644511149
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2098_
timestamp 1644511149
transform -1 0 22264 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2099_
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _2100_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2101_
timestamp 1644511149
transform -1 0 17296 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2102_
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2103_
timestamp 1644511149
transform -1 0 9844 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2104_
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _2105_
timestamp 1644511149
transform -1 0 8096 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2106_
timestamp 1644511149
transform 1 0 9200 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2107_
timestamp 1644511149
transform 1 0 11868 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2108_
timestamp 1644511149
transform -1 0 15824 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2109_
timestamp 1644511149
transform -1 0 15088 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _2110_
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2111_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _2112_
timestamp 1644511149
transform -1 0 10948 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _2113_
timestamp 1644511149
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _2114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19872 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2115_
timestamp 1644511149
transform -1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2116_
timestamp 1644511149
transform 1 0 10764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2117_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2118_
timestamp 1644511149
transform 1 0 14720 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2119_
timestamp 1644511149
transform 1 0 11224 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_1  _2120_
timestamp 1644511149
transform 1 0 10304 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2121_
timestamp 1644511149
transform -1 0 9844 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2122_
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2123_
timestamp 1644511149
transform -1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2124_
timestamp 1644511149
transform -1 0 19504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2125_
timestamp 1644511149
transform -1 0 18308 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2126_
timestamp 1644511149
transform -1 0 10488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2127_
timestamp 1644511149
transform 1 0 9384 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2128_
timestamp 1644511149
transform -1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2129_
timestamp 1644511149
transform 1 0 30728 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2130_
timestamp 1644511149
transform -1 0 32016 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2131_
timestamp 1644511149
transform -1 0 32660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2132_
timestamp 1644511149
transform 1 0 33028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2133_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2134_
timestamp 1644511149
transform 1 0 35328 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2135_
timestamp 1644511149
transform 1 0 31372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2136_
timestamp 1644511149
transform 1 0 35512 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2137_
timestamp 1644511149
transform 1 0 36432 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2138_
timestamp 1644511149
transform 1 0 35236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2139_
timestamp 1644511149
transform -1 0 34684 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2140_
timestamp 1644511149
transform -1 0 30636 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2141_
timestamp 1644511149
transform -1 0 23920 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _2142_
timestamp 1644511149
transform 1 0 26036 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2143_
timestamp 1644511149
transform 1 0 29716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2144_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2145_
timestamp 1644511149
transform -1 0 26220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2146_
timestamp 1644511149
transform 1 0 30084 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2147_
timestamp 1644511149
transform 1 0 29808 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2148_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2149_
timestamp 1644511149
transform -1 0 33396 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2150_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2151_
timestamp 1644511149
transform -1 0 32384 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2152_
timestamp 1644511149
transform -1 0 30728 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2153_
timestamp 1644511149
transform -1 0 25300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2154_
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2155_
timestamp 1644511149
transform 1 0 22632 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2156_
timestamp 1644511149
transform -1 0 22448 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2157_
timestamp 1644511149
transform -1 0 23276 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2158_
timestamp 1644511149
transform 1 0 23828 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2159_
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2160_
timestamp 1644511149
transform -1 0 24748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2161_
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2162_
timestamp 1644511149
transform -1 0 22632 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2163_
timestamp 1644511149
transform -1 0 27508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2164_
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2165_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2166_
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2167_
timestamp 1644511149
transform 1 0 24748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2168_
timestamp 1644511149
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2169_
timestamp 1644511149
transform -1 0 17204 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2170_
timestamp 1644511149
transform -1 0 19504 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2171_
timestamp 1644511149
transform -1 0 19964 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2172_
timestamp 1644511149
transform -1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2173_
timestamp 1644511149
transform -1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2174_
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2175_
timestamp 1644511149
transform 1 0 12144 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2176_
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2177_
timestamp 1644511149
transform -1 0 10028 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2178_
timestamp 1644511149
transform -1 0 10948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2179_
timestamp 1644511149
transform -1 0 9016 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2180_
timestamp 1644511149
transform 1 0 9016 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2181_
timestamp 1644511149
transform 1 0 8372 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2182_
timestamp 1644511149
transform -1 0 5888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2183_
timestamp 1644511149
transform -1 0 5244 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2184_
timestamp 1644511149
transform -1 0 4968 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2185_
timestamp 1644511149
transform -1 0 10856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2186_
timestamp 1644511149
transform -1 0 6716 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2187_
timestamp 1644511149
transform -1 0 10304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2188_
timestamp 1644511149
transform 1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2189_
timestamp 1644511149
transform 1 0 10120 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2190_
timestamp 1644511149
transform 1 0 8464 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2191_
timestamp 1644511149
transform 1 0 13524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2192_
timestamp 1644511149
transform -1 0 14996 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2193_
timestamp 1644511149
transform -1 0 14536 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2194_
timestamp 1644511149
transform 1 0 20148 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2195_
timestamp 1644511149
transform -1 0 16008 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2196_
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2197_
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2198_
timestamp 1644511149
transform 1 0 17296 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2199_
timestamp 1644511149
transform -1 0 15180 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2200_
timestamp 1644511149
transform 1 0 21712 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2201_
timestamp 1644511149
transform -1 0 21068 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2202_
timestamp 1644511149
transform 1 0 17020 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2203_
timestamp 1644511149
transform 1 0 23184 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2204_
timestamp 1644511149
transform -1 0 24748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2205_
timestamp 1644511149
transform -1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2206_
timestamp 1644511149
transform -1 0 20792 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2207_
timestamp 1644511149
transform -1 0 20884 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2208_
timestamp 1644511149
transform -1 0 20148 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2209_
timestamp 1644511149
transform -1 0 22816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2210_
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2211_
timestamp 1644511149
transform -1 0 25668 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2212_
timestamp 1644511149
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2213_
timestamp 1644511149
transform -1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2214_
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2215_
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2216_
timestamp 1644511149
transform 1 0 30544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2217_
timestamp 1644511149
transform -1 0 30176 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2218_
timestamp 1644511149
transform -1 0 30084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2219_
timestamp 1644511149
transform -1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2220_
timestamp 1644511149
transform -1 0 33028 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2221_
timestamp 1644511149
transform 1 0 33396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2222_
timestamp 1644511149
transform 1 0 35236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2223_
timestamp 1644511149
transform 1 0 35512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2224_
timestamp 1644511149
transform 1 0 34132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2225_
timestamp 1644511149
transform -1 0 33580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2226_
timestamp 1644511149
transform -1 0 35604 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2227_
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2228_
timestamp 1644511149
transform 1 0 36432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2229_
timestamp 1644511149
transform -1 0 36708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2230_
timestamp 1644511149
transform -1 0 35880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2231_
timestamp 1644511149
transform -1 0 35052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2232_
timestamp 1644511149
transform -1 0 35880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2233_
timestamp 1644511149
transform 1 0 34960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2234_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2235_
timestamp 1644511149
transform 1 0 30360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2236_
timestamp 1644511149
transform 1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2237_
timestamp 1644511149
transform 1 0 35512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2238_
timestamp 1644511149
transform 1 0 32936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2239_
timestamp 1644511149
transform 1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2240_
timestamp 1644511149
transform -1 0 29808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2241_
timestamp 1644511149
transform 1 0 26864 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2242_
timestamp 1644511149
transform 1 0 24840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2243_
timestamp 1644511149
transform 1 0 27416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2244_
timestamp 1644511149
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2245_
timestamp 1644511149
transform 1 0 24932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2246_
timestamp 1644511149
transform -1 0 23920 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2247_
timestamp 1644511149
transform -1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2248_
timestamp 1644511149
transform -1 0 23920 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2249_
timestamp 1644511149
transform 1 0 22356 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2250_
timestamp 1644511149
transform 1 0 21712 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2251_
timestamp 1644511149
transform -1 0 21344 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2252_
timestamp 1644511149
transform -1 0 20700 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2253_
timestamp 1644511149
transform 1 0 27600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2254_
timestamp 1644511149
transform -1 0 26956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2255_
timestamp 1644511149
transform -1 0 21344 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2256_
timestamp 1644511149
transform 1 0 27232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2257_
timestamp 1644511149
transform -1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2258_
timestamp 1644511149
transform 1 0 32108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2259_
timestamp 1644511149
transform -1 0 29900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2260_
timestamp 1644511149
transform -1 0 30728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2261_
timestamp 1644511149
transform -1 0 31096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2262_
timestamp 1644511149
transform 1 0 31096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2263_
timestamp 1644511149
transform -1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2264_
timestamp 1644511149
transform -1 0 27876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2265_
timestamp 1644511149
transform -1 0 22172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2266_
timestamp 1644511149
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2267_
timestamp 1644511149
transform 1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2268_
timestamp 1644511149
transform -1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2269_
timestamp 1644511149
transform -1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2270_
timestamp 1644511149
transform -1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2271_
timestamp 1644511149
transform -1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2272_
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2273_
timestamp 1644511149
transform 1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2274_
timestamp 1644511149
transform -1 0 15640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2275_
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2276_
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2277_
timestamp 1644511149
transform -1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2278_
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2279_
timestamp 1644511149
transform -1 0 14996 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2280_
timestamp 1644511149
transform -1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2281_
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2282_
timestamp 1644511149
transform -1 0 14168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2283_
timestamp 1644511149
transform 1 0 15640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2284_
timestamp 1644511149
transform -1 0 12788 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2285_
timestamp 1644511149
transform 1 0 14352 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2286_
timestamp 1644511149
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2287_
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2288_
timestamp 1644511149
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2289_
timestamp 1644511149
transform -1 0 26312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2290_
timestamp 1644511149
transform -1 0 19596 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2291_
timestamp 1644511149
transform 1 0 13984 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2292_
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _2293_
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2294_
timestamp 1644511149
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2295_
timestamp 1644511149
transform 1 0 8648 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2296_
timestamp 1644511149
transform 1 0 6808 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _2297_
timestamp 1644511149
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2298_
timestamp 1644511149
transform -1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2299_
timestamp 1644511149
transform -1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2300_
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _2301_
timestamp 1644511149
transform 1 0 5060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2302_
timestamp 1644511149
transform -1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2303_
timestamp 1644511149
transform -1 0 9476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2304_
timestamp 1644511149
transform 1 0 7636 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2305_
timestamp 1644511149
transform 1 0 7452 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _2306_
timestamp 1644511149
transform -1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2307_
timestamp 1644511149
transform -1 0 6440 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2308_
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _2309_
timestamp 1644511149
transform 1 0 8648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2310_
timestamp 1644511149
transform -1 0 7084 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2311_
timestamp 1644511149
transform -1 0 7084 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2312_
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2313_
timestamp 1644511149
transform -1 0 9200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2314_
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2315_
timestamp 1644511149
transform -1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2316_
timestamp 1644511149
transform -1 0 8832 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2317_
timestamp 1644511149
transform 1 0 8280 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2318_
timestamp 1644511149
transform -1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2319_
timestamp 1644511149
transform 1 0 7636 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2320_
timestamp 1644511149
transform -1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2321_
timestamp 1644511149
transform 1 0 7544 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2322_
timestamp 1644511149
transform -1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _2323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20056 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2324_
timestamp 1644511149
transform -1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2325_
timestamp 1644511149
transform -1 0 14812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2326_
timestamp 1644511149
transform 1 0 9476 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2327_
timestamp 1644511149
transform -1 0 9936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2328_
timestamp 1644511149
transform 1 0 10396 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2329_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _2330_
timestamp 1644511149
transform 1 0 9844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2331_
timestamp 1644511149
transform -1 0 12052 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2332_
timestamp 1644511149
transform 1 0 10488 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2333_
timestamp 1644511149
transform -1 0 12880 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2334_
timestamp 1644511149
transform -1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _2335_
timestamp 1644511149
transform 1 0 11040 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2336_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2337_
timestamp 1644511149
transform -1 0 12880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2338_
timestamp 1644511149
transform 1 0 12512 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2339_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2340_
timestamp 1644511149
transform 1 0 11868 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2341_
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2342_
timestamp 1644511149
transform 1 0 11960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2343_
timestamp 1644511149
transform 1 0 13524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2344_
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2345_
timestamp 1644511149
transform -1 0 14352 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2346_
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2347_
timestamp 1644511149
transform 1 0 16928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2348_
timestamp 1644511149
transform 1 0 16836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2349_
timestamp 1644511149
transform -1 0 16928 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2350_
timestamp 1644511149
transform -1 0 16376 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2351_
timestamp 1644511149
transform 1 0 15088 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2352_
timestamp 1644511149
transform -1 0 13708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2353_
timestamp 1644511149
transform -1 0 16192 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2354_
timestamp 1644511149
transform -1 0 15548 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2355_
timestamp 1644511149
transform 1 0 14720 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2356_
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2357_
timestamp 1644511149
transform 1 0 14352 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2358_
timestamp 1644511149
transform -1 0 15640 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2359_
timestamp 1644511149
transform 1 0 14628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2360_
timestamp 1644511149
transform -1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2361_
timestamp 1644511149
transform -1 0 14812 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2362_
timestamp 1644511149
transform 1 0 16468 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _2363_
timestamp 1644511149
transform -1 0 17020 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2364_
timestamp 1644511149
transform -1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2365_
timestamp 1644511149
transform 1 0 17940 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2366_
timestamp 1644511149
transform -1 0 16008 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2367_
timestamp 1644511149
transform -1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2368_
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2369_
timestamp 1644511149
transform -1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2370_
timestamp 1644511149
transform 1 0 15364 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2371_
timestamp 1644511149
transform 1 0 15180 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2372_
timestamp 1644511149
transform -1 0 17296 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2373_
timestamp 1644511149
transform -1 0 17020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2374_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2375_
timestamp 1644511149
transform -1 0 18216 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2376_
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2377_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2378_
timestamp 1644511149
transform -1 0 20424 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2379_
timestamp 1644511149
transform 1 0 18492 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2380_
timestamp 1644511149
transform -1 0 18124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2381_
timestamp 1644511149
transform 1 0 15732 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _2382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _2383_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2384_
timestamp 1644511149
transform -1 0 20608 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2385_
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2386_
timestamp 1644511149
transform -1 0 16192 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2387_
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2388_
timestamp 1644511149
transform -1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2389_
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2390_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2391_
timestamp 1644511149
transform -1 0 13340 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2392_
timestamp 1644511149
transform -1 0 11040 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2393_
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2394_
timestamp 1644511149
transform -1 0 13524 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2395_
timestamp 1644511149
transform 1 0 12972 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2396_
timestamp 1644511149
transform -1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2397_
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2398_
timestamp 1644511149
transform -1 0 14720 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2399_
timestamp 1644511149
transform -1 0 13248 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2400_
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2401_
timestamp 1644511149
transform -1 0 11040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2402_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2403_
timestamp 1644511149
transform 1 0 11408 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2404_
timestamp 1644511149
transform 1 0 10212 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2405_
timestamp 1644511149
transform -1 0 10028 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2406_
timestamp 1644511149
transform 1 0 9200 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2407_
timestamp 1644511149
transform 1 0 12512 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2408_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2409_
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2410_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8004 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2411_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2413_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2414_
timestamp 1644511149
transform 1 0 30268 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2415_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2416_
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2417_
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2418_
timestamp 1644511149
transform 1 0 34500 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2419_
timestamp 1644511149
transform 1 0 34592 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2420_
timestamp 1644511149
transform 1 0 34224 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2421_
timestamp 1644511149
transform -1 0 33856 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2422_
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2423_
timestamp 1644511149
transform -1 0 31004 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2424_
timestamp 1644511149
transform 1 0 26036 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2425_
timestamp 1644511149
transform 1 0 24840 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2426_
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2427_
timestamp 1644511149
transform -1 0 31372 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2428_
timestamp 1644511149
transform 1 0 32016 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2429_
timestamp 1644511149
transform 1 0 33396 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2430_
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2431_
timestamp 1644511149
transform -1 0 30820 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2432_
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2433_
timestamp 1644511149
transform 1 0 21620 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2434_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2435_
timestamp 1644511149
transform 1 0 21896 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2436_
timestamp 1644511149
transform -1 0 27232 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2437_
timestamp 1644511149
transform -1 0 26312 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2438_
timestamp 1644511149
transform -1 0 25208 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2439_
timestamp 1644511149
transform -1 0 26220 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2440_
timestamp 1644511149
transform 1 0 26128 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2441_
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2442_
timestamp 1644511149
transform 1 0 27048 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2443_
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2444_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2445_
timestamp 1644511149
transform 1 0 15364 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2446_
timestamp 1644511149
transform 1 0 17020 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2447_
timestamp 1644511149
transform 1 0 15456 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2448_
timestamp 1644511149
transform -1 0 15916 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2449_
timestamp 1644511149
transform 1 0 11684 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2450_
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2451_
timestamp 1644511149
transform 1 0 8464 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2452_
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2453_
timestamp 1644511149
transform -1 0 10764 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2454_
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2455_
timestamp 1644511149
transform -1 0 6624 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2456_
timestamp 1644511149
transform -1 0 6164 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2457_
timestamp 1644511149
transform -1 0 6256 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2458_
timestamp 1644511149
transform -1 0 6900 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2459_
timestamp 1644511149
transform -1 0 10672 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2460_
timestamp 1644511149
transform 1 0 6440 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2461_
timestamp 1644511149
transform 1 0 9108 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2462_
timestamp 1644511149
transform -1 0 10764 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2463_
timestamp 1644511149
transform -1 0 13616 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2464_
timestamp 1644511149
transform 1 0 12328 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2465_
timestamp 1644511149
transform 1 0 14444 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2466_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2467_
timestamp 1644511149
transform 1 0 13248 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2468_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2469_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2470_
timestamp 1644511149
transform -1 0 21344 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2471_
timestamp 1644511149
transform -1 0 21160 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2472_
timestamp 1644511149
transform -1 0 19504 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2473_
timestamp 1644511149
transform 1 0 19688 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2474_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2475_
timestamp 1644511149
transform -1 0 21344 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2476_
timestamp 1644511149
transform -1 0 21068 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2477_
timestamp 1644511149
transform 1 0 20792 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2478_
timestamp 1644511149
transform 1 0 23736 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2479_
timestamp 1644511149
transform 1 0 23368 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2480_
timestamp 1644511149
transform -1 0 26220 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2481_
timestamp 1644511149
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2482_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2483_
timestamp 1644511149
transform 1 0 28244 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2484_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2485_
timestamp 1644511149
transform 1 0 30452 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2486_
timestamp 1644511149
transform -1 0 32752 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2487_
timestamp 1644511149
transform 1 0 32016 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2488_
timestamp 1644511149
transform 1 0 34960 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2489_
timestamp 1644511149
transform -1 0 36800 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2490_
timestamp 1644511149
transform 1 0 34776 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2491_
timestamp 1644511149
transform 1 0 33948 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2492_
timestamp 1644511149
transform -1 0 37996 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2493_
timestamp 1644511149
transform 1 0 34224 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2494_
timestamp 1644511149
transform -1 0 36616 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2495_
timestamp 1644511149
transform 1 0 33028 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2496_
timestamp 1644511149
transform 1 0 32384 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2497_
timestamp 1644511149
transform -1 0 36800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2498_
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2499_
timestamp 1644511149
transform 1 0 32384 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2500_
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2501_
timestamp 1644511149
transform -1 0 32016 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2502_
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2503_
timestamp 1644511149
transform -1 0 30268 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2504_
timestamp 1644511149
transform 1 0 27048 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2505_
timestamp 1644511149
transform 1 0 27876 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2506_
timestamp 1644511149
transform -1 0 31464 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2507_
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2508_
timestamp 1644511149
transform -1 0 24932 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2509_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2510_
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2511_
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2512_
timestamp 1644511149
transform 1 0 19964 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2513_
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2514_
timestamp 1644511149
transform -1 0 26220 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2515_
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2516_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2517_
timestamp 1644511149
transform 1 0 22816 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2518_
timestamp 1644511149
transform 1 0 24932 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2519_
timestamp 1644511149
transform 1 0 28704 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2520_
timestamp 1644511149
transform 1 0 28612 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2521_
timestamp 1644511149
transform 1 0 28244 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2522_
timestamp 1644511149
transform -1 0 28888 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2523_
timestamp 1644511149
transform -1 0 26496 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2524_
timestamp 1644511149
transform -1 0 26864 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2525_
timestamp 1644511149
transform -1 0 24840 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2526_
timestamp 1644511149
transform 1 0 21804 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2527_
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2528_
timestamp 1644511149
transform 1 0 19412 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2529_
timestamp 1644511149
transform 1 0 15272 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2530_
timestamp 1644511149
transform 1 0 14536 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2531_
timestamp 1644511149
transform 1 0 16836 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2532_
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2533_
timestamp 1644511149
transform 1 0 13064 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2534_
timestamp 1644511149
transform -1 0 15916 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2535_
timestamp 1644511149
transform 1 0 12880 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2536_
timestamp 1644511149
transform -1 0 16744 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2537_
timestamp 1644511149
transform -1 0 16008 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2538_
timestamp 1644511149
transform -1 0 16468 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2539_
timestamp 1644511149
transform 1 0 13892 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2540_
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2541_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2542_
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2543_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2544_
timestamp 1644511149
transform -1 0 23000 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2545_
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2546_
timestamp 1644511149
transform 1 0 4416 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2547_
timestamp 1644511149
transform 1 0 4324 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2548_
timestamp 1644511149
transform 1 0 4324 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2549_
timestamp 1644511149
transform 1 0 5244 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2550_
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2551_
timestamp 1644511149
transform 1 0 6624 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2552_
timestamp 1644511149
transform 1 0 9568 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2553_
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2554_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2555_
timestamp 1644511149
transform 1 0 10580 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2556_
timestamp 1644511149
transform 1 0 11684 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2557_
timestamp 1644511149
transform 1 0 12788 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2558_
timestamp 1644511149
transform -1 0 18768 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2559_
timestamp 1644511149
transform -1 0 17388 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2560_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2561_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2562_
timestamp 1644511149
transform -1 0 18124 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2563_
timestamp 1644511149
transform 1 0 14720 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2564_
timestamp 1644511149
transform -1 0 18124 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2565_
timestamp 1644511149
transform -1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2566_
timestamp 1644511149
transform -1 0 21436 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2567_
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2568_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2569_
timestamp 1644511149
transform 1 0 12420 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2570_
timestamp 1644511149
transform 1 0 12144 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2571_
timestamp 1644511149
transform 1 0 13616 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2572_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2573_
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2574_
timestamp 1644511149
transform 1 0 7728 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _2575__3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2576__4
timestamp 1644511149
transform 1 0 1472 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2577__5
timestamp 1644511149
transform -1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2578__6
timestamp 1644511149
transform -1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2579__7
timestamp 1644511149
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2580__8
timestamp 1644511149
transform 1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2581__9
timestamp 1644511149
transform 1 0 33672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2582__10
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2583__11
timestamp 1644511149
transform 1 0 35880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2584__12
timestamp 1644511149
transform -1 0 36800 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2585__13
timestamp 1644511149
transform 1 0 37628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2586__14
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2587__15
timestamp 1644511149
transform 1 0 35604 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2588__16
timestamp 1644511149
transform -1 0 8004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2589__17
timestamp 1644511149
transform 1 0 23460 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2590__18
timestamp 1644511149
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2591__19
timestamp 1644511149
transform 1 0 35604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2592__20
timestamp 1644511149
transform 1 0 37628 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2593__21
timestamp 1644511149
transform -1 0 8004 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2594__22
timestamp 1644511149
transform 1 0 37628 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2595__23
timestamp 1644511149
transform 1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2596__24
timestamp 1644511149
transform 1 0 37904 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2597__25
timestamp 1644511149
transform -1 0 24656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2598__26
timestamp 1644511149
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2599__27
timestamp 1644511149
transform 1 0 34960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2600__28
timestamp 1644511149
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2601__29
timestamp 1644511149
transform -1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2602__30
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2603__31
timestamp 1644511149
transform -1 0 35236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2604__32
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2605__33
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2606__34
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2607__35
timestamp 1644511149
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2608__36
timestamp 1644511149
transform 1 0 25208 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2609__37
timestamp 1644511149
transform -1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2610__38
timestamp 1644511149
transform -1 0 3864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2611__39
timestamp 1644511149
transform -1 0 36800 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2612__40
timestamp 1644511149
transform -1 0 17940 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2613__41
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2614__42
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2615__43
timestamp 1644511149
transform -1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2616__44
timestamp 1644511149
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2617__45
timestamp 1644511149
transform 1 0 37904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2618__46
timestamp 1644511149
transform -1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2619__47
timestamp 1644511149
transform 1 0 1472 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2620__48
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2621__49
timestamp 1644511149
transform 1 0 35236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2622__50
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2623__51
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2624__52
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2625__53
timestamp 1644511149
transform -1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2626__54
timestamp 1644511149
transform 1 0 37628 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2627__55
timestamp 1644511149
transform -1 0 22724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2628__56
timestamp 1644511149
transform -1 0 30452 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2629__57
timestamp 1644511149
transform -1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2630__58
timestamp 1644511149
transform -1 0 32384 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2631__59
timestamp 1644511149
transform 1 0 13064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2632__60
timestamp 1644511149
transform 1 0 37904 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2633__61
timestamp 1644511149
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2634__62
timestamp 1644511149
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2635__63
timestamp 1644511149
transform 1 0 2392 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2636__64
timestamp 1644511149
transform -1 0 37904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2637__65
timestamp 1644511149
transform -1 0 36800 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2638__66
timestamp 1644511149
transform 1 0 35236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2639__67
timestamp 1644511149
transform 1 0 14720 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2640__68
timestamp 1644511149
transform 1 0 35604 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2641__69
timestamp 1644511149
transform -1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2642__70
timestamp 1644511149
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2643__71
timestamp 1644511149
transform -1 0 32660 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2644__72
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2645__73
timestamp 1644511149
transform 1 0 35880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2646__74
timestamp 1644511149
transform -1 0 2208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2647__75
timestamp 1644511149
transform 1 0 37904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2648__76
timestamp 1644511149
transform -1 0 10028 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2649__77
timestamp 1644511149
transform -1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2650__78
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2651__79
timestamp 1644511149
transform -1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2652__80
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2653__81
timestamp 1644511149
transform 1 0 33948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2654__82
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2655__83
timestamp 1644511149
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2656__84
timestamp 1644511149
transform 1 0 10396 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2657__85
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2658__86
timestamp 1644511149
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2659__87
timestamp 1644511149
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2660__88
timestamp 1644511149
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2661__89
timestamp 1644511149
transform 1 0 32660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2662__90
timestamp 1644511149
transform 1 0 1932 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2663__91
timestamp 1644511149
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2664__92
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2665__93
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2666__94
timestamp 1644511149
transform -1 0 35880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2667__95
timestamp 1644511149
transform 1 0 35880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2668__96
timestamp 1644511149
transform -1 0 23276 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2669__97
timestamp 1644511149
transform -1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2670__98
timestamp 1644511149
transform -1 0 37260 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2671__99
timestamp 1644511149
transform 1 0 3036 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2672__100
timestamp 1644511149
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2673__101
timestamp 1644511149
transform -1 0 1840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2674__102
timestamp 1644511149
transform -1 0 35880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2675__103
timestamp 1644511149
transform -1 0 8648 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2676__104
timestamp 1644511149
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2677__105
timestamp 1644511149
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2678__106
timestamp 1644511149
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2679_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2680_
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2681_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2682_
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2683_
timestamp 1644511149
transform 1 0 35420 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2684_
timestamp 1644511149
transform -1 0 4416 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2685_
timestamp 1644511149
transform 1 0 36248 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2686_
timestamp 1644511149
transform -1 0 3312 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2687_
timestamp 1644511149
transform 1 0 36248 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2688_
timestamp 1644511149
transform 1 0 36248 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2689_
timestamp 1644511149
transform -1 0 38180 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2690_
timestamp 1644511149
transform 1 0 18952 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2691_
timestamp 1644511149
transform 1 0 36248 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2692_
timestamp 1644511149
transform -1 0 5796 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2693_
timestamp 1644511149
transform -1 0 23736 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2694_
timestamp 1644511149
transform -1 0 4600 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2695_
timestamp 1644511149
transform 1 0 36248 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2696_
timestamp 1644511149
transform -1 0 38180 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2697_
timestamp 1644511149
transform -1 0 5888 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2698_
timestamp 1644511149
transform -1 0 38180 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2699_
timestamp 1644511149
transform -1 0 5888 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2700_
timestamp 1644511149
transform -1 0 38180 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2701_
timestamp 1644511149
transform 1 0 24104 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2702_
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2703_
timestamp 1644511149
transform 1 0 36248 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2704_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2705_
timestamp 1644511149
transform 1 0 35696 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2706_
timestamp 1644511149
transform -1 0 3312 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2707_
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2708_
timestamp 1644511149
transform -1 0 5980 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2709_
timestamp 1644511149
transform 1 0 36248 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2710_
timestamp 1644511149
transform 1 0 34868 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2711_
timestamp 1644511149
transform 1 0 34868 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2712_
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2713_
timestamp 1644511149
transform 1 0 4968 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2714_
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2715_
timestamp 1644511149
transform 1 0 36248 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2716_
timestamp 1644511149
transform 1 0 17664 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2717_
timestamp 1644511149
transform 1 0 34868 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2718_
timestamp 1644511149
transform -1 0 3312 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2719_
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2720_
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2721_
timestamp 1644511149
transform -1 0 38180 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2722_
timestamp 1644511149
transform -1 0 3312 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2723_
timestamp 1644511149
transform 1 0 1656 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2724_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2725_
timestamp 1644511149
transform 1 0 36248 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2726_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2727_
timestamp 1644511149
transform 1 0 36248 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2728_
timestamp 1644511149
transform 1 0 36156 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2729_
timestamp 1644511149
transform 1 0 36248 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2730_
timestamp 1644511149
transform 1 0 1656 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2731_
timestamp 1644511149
transform 1 0 31648 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2732_
timestamp 1644511149
transform -1 0 3312 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2733_
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2734_
timestamp 1644511149
transform -1 0 38180 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2735_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2736_
timestamp 1644511149
transform 1 0 29072 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2737_
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2738_
timestamp 1644511149
transform 1 0 29716 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2739_
timestamp 1644511149
transform -1 0 13892 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2740_
timestamp 1644511149
transform -1 0 38180 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2741_
timestamp 1644511149
transform -1 0 3680 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2742_
timestamp 1644511149
transform 1 0 1564 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2743_
timestamp 1644511149
transform -1 0 3496 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2744_
timestamp 1644511149
transform 1 0 36248 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2745_
timestamp 1644511149
transform 1 0 36248 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2746_
timestamp 1644511149
transform 1 0 36248 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2747_
timestamp 1644511149
transform -1 0 16192 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2748_
timestamp 1644511149
transform -1 0 36800 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2749_
timestamp 1644511149
transform -1 0 22632 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2750_
timestamp 1644511149
transform 1 0 31004 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2751_
timestamp 1644511149
transform 1 0 32384 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2752_
timestamp 1644511149
transform 1 0 19320 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2753_
timestamp 1644511149
transform -1 0 36800 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2754_
timestamp 1644511149
transform 1 0 1840 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2755_
timestamp 1644511149
transform -1 0 38180 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2756_
timestamp 1644511149
transform 1 0 9752 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2757_
timestamp 1644511149
transform -1 0 5704 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2758_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2759_
timestamp 1644511149
transform 1 0 1840 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2760_
timestamp 1644511149
transform 1 0 34868 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2761_
timestamp 1644511149
transform 1 0 36248 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2762_
timestamp 1644511149
transform -1 0 36800 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2763_
timestamp 1644511149
transform -1 0 10856 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2764_
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2765_
timestamp 1644511149
transform -1 0 36800 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2766_
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2767_
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2768_
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2769_
timestamp 1644511149
transform 1 0 34868 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2770_
timestamp 1644511149
transform -1 0 3312 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2771_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2772_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2773_
timestamp 1644511149
transform 1 0 19412 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2774_
timestamp 1644511149
transform -1 0 34224 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2775_
timestamp 1644511149
transform 1 0 36248 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2776_
timestamp 1644511149
transform 1 0 22632 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2777_
timestamp 1644511149
transform 1 0 32568 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2778_
timestamp 1644511149
transform 1 0 36248 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2779_
timestamp 1644511149
transform -1 0 5704 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2780_
timestamp 1644511149
transform 1 0 32200 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2781_
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2782_
timestamp 1644511149
transform 1 0 35604 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2783_
timestamp 1644511149
transform 1 0 8372 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2784_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2785_
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2786_
timestamp 1644511149
transform -1 0 3312 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22448 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform -1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 16192 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 28980 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform -1 0 30912 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 12972 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 14904 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 16928 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform -1 0 27324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 28704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 25392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1644511149
transform -1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1644511149
transform -1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1644511149
transform -1 0 11868 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1644511149
transform -1 0 17572 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1644511149
transform -1 0 26312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1644511149
transform -1 0 25852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1644511149
transform -1 0 31464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1644511149
transform 1 0 31280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1644511149
transform 1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1644511149
transform -1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1644511149
transform 1 0 33856 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1644511149
transform -1 0 31648 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform -1 0 38180 0 -1 6528
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 36668 800 36908 6 active
port 0 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 21886 39200 21998 40000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s -10 39200 102 40000 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 39200 33268 40000 33508 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 14802 39200 14914 40000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 39200 35308 40000 35548 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 39200 3348 40000 3588 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 7718 39200 7830 40000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 9650 39200 9762 40000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 39200 12868 40000 13108 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 7074 39200 7186 40000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 5142 39200 5254 40000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 39200 8788 40000 9028 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 39274 39200 39386 40000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 39200 15588 40000 15828 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 30258 39200 30370 40000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 34766 39200 34878 40000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 39200 25108 40000 25348 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 35410 39200 35522 40000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 22530 39200 22642 40000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 39200 24428 40000 24668 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 39200 38028 40000 38268 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 39200 26468 40000 26708 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 6430 39200 6542 40000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 io_oeb[0]
port 39 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 io_oeb[10]
port 40 nsew signal bidirectional
rlabel metal3 s 39200 22388 40000 22628 6 io_oeb[11]
port 41 nsew signal bidirectional
rlabel metal3 s 39200 11508 40000 11748 6 io_oeb[12]
port 42 nsew signal bidirectional
rlabel metal3 s 39200 10828 40000 11068 6 io_oeb[13]
port 43 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 44 nsew signal bidirectional
rlabel metal2 s 10938 39200 11050 40000 6 io_oeb[15]
port 45 nsew signal bidirectional
rlabel metal3 s 39200 1988 40000 2228 6 io_oeb[16]
port 46 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 io_oeb[17]
port 47 nsew signal bidirectional
rlabel metal2 s 28326 39200 28438 40000 6 io_oeb[18]
port 48 nsew signal bidirectional
rlabel metal2 s 11582 39200 11694 40000 6 io_oeb[19]
port 49 nsew signal bidirectional
rlabel metal2 s 31546 0 31658 800 6 io_oeb[1]
port 50 nsew signal bidirectional
rlabel metal3 s 39200 16948 40000 17188 6 io_oeb[20]
port 51 nsew signal bidirectional
rlabel metal2 s 1278 39200 1390 40000 6 io_oeb[21]
port 52 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 53 nsew signal bidirectional
rlabel metal2 s 19954 39200 20066 40000 6 io_oeb[23]
port 54 nsew signal bidirectional
rlabel metal2 s 20598 39200 20710 40000 6 io_oeb[24]
port 55 nsew signal bidirectional
rlabel metal2 s 37986 0 38098 800 6 io_oeb[25]
port 56 nsew signal bidirectional
rlabel metal3 s 39200 31228 40000 31468 6 io_oeb[26]
port 57 nsew signal bidirectional
rlabel metal2 s 23174 39200 23286 40000 6 io_oeb[27]
port 58 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 io_oeb[28]
port 59 nsew signal bidirectional
rlabel metal3 s 39200 25788 40000 26028 6 io_oeb[29]
port 60 nsew signal bidirectional
rlabel metal2 s 32834 39200 32946 40000 6 io_oeb[2]
port 61 nsew signal bidirectional
rlabel metal2 s 1922 39200 2034 40000 6 io_oeb[30]
port 62 nsew signal bidirectional
rlabel metal2 s 32834 0 32946 800 6 io_oeb[31]
port 63 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 io_oeb[32]
port 64 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 io_oeb[33]
port 65 nsew signal bidirectional
rlabel metal2 s 9006 39200 9118 40000 6 io_oeb[34]
port 66 nsew signal bidirectional
rlabel metal3 s 0 17628 800 17868 6 io_oeb[35]
port 67 nsew signal bidirectional
rlabel metal3 s 0 8788 800 9028 6 io_oeb[36]
port 68 nsew signal bidirectional
rlabel metal3 s 0 14228 800 14468 6 io_oeb[37]
port 69 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 io_oeb[3]
port 70 nsew signal bidirectional
rlabel metal3 s 39200 -52 40000 188 6 io_oeb[4]
port 71 nsew signal bidirectional
rlabel metal3 s 0 25788 800 26028 6 io_oeb[5]
port 72 nsew signal bidirectional
rlabel metal3 s 39200 14228 40000 14468 6 io_oeb[6]
port 73 nsew signal bidirectional
rlabel metal2 s 10294 39200 10406 40000 6 io_oeb[7]
port 74 nsew signal bidirectional
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 75 nsew signal bidirectional
rlabel metal2 s 8362 0 8474 800 6 io_oeb[9]
port 76 nsew signal bidirectional
rlabel metal3 s 39200 37348 40000 37588 6 io_out[0]
port 77 nsew signal bidirectional
rlabel metal3 s 39200 21708 40000 21948 6 io_out[10]
port 78 nsew signal bidirectional
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal bidirectional
rlabel metal3 s 0 6068 800 6308 6 io_out[12]
port 80 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 io_out[13]
port 81 nsew signal bidirectional
rlabel metal3 s 39200 31908 40000 32148 6 io_out[14]
port 82 nsew signal bidirectional
rlabel metal3 s 0 33268 800 33508 6 io_out[15]
port 83 nsew signal bidirectional
rlabel metal3 s 39200 21028 40000 21268 6 io_out[16]
port 84 nsew signal bidirectional
rlabel metal2 s 36698 39200 36810 40000 6 io_out[17]
port 85 nsew signal bidirectional
rlabel metal2 s 37342 0 37454 800 6 io_out[18]
port 86 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 io_out[19]
port 87 nsew signal bidirectional
rlabel metal2 s 26394 39200 26506 40000 6 io_out[1]
port 88 nsew signal bidirectional
rlabel metal2 s 32190 39200 32302 40000 6 io_out[20]
port 89 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 io_out[21]
port 90 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 io_out[22]
port 91 nsew signal bidirectional
rlabel metal3 s 39200 18308 40000 18548 6 io_out[23]
port 92 nsew signal bidirectional
rlabel metal2 s 21886 0 21998 800 6 io_out[24]
port 93 nsew signal bidirectional
rlabel metal2 s 29614 39200 29726 40000 6 io_out[25]
port 94 nsew signal bidirectional
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 95 nsew signal bidirectional
rlabel metal2 s 30902 39200 31014 40000 6 io_out[27]
port 96 nsew signal bidirectional
rlabel metal2 s 13514 0 13626 800 6 io_out[28]
port 97 nsew signal bidirectional
rlabel metal3 s 39200 628 40000 868 6 io_out[29]
port 98 nsew signal bidirectional
rlabel metal2 s 5786 0 5898 800 6 io_out[2]
port 99 nsew signal bidirectional
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 100 nsew signal bidirectional
rlabel metal3 s 0 11508 800 11748 6 io_out[31]
port 101 nsew signal bidirectional
rlabel metal3 s 0 37348 800 37588 6 io_out[32]
port 102 nsew signal bidirectional
rlabel metal3 s 39200 5388 40000 5628 6 io_out[33]
port 103 nsew signal bidirectional
rlabel metal3 s 39200 32588 40000 32828 6 io_out[34]
port 104 nsew signal bidirectional
rlabel metal3 s 39200 30548 40000 30788 6 io_out[35]
port 105 nsew signal bidirectional
rlabel metal2 s 12226 39200 12338 40000 6 io_out[36]
port 106 nsew signal bidirectional
rlabel metal3 s 39200 35988 40000 36228 6 io_out[37]
port 107 nsew signal bidirectional
rlabel metal3 s 0 34628 800 34868 6 io_out[3]
port 108 nsew signal bidirectional
rlabel metal3 s 39200 23748 40000 23988 6 io_out[4]
port 109 nsew signal bidirectional
rlabel metal2 s 18022 39200 18134 40000 6 io_out[5]
port 110 nsew signal bidirectional
rlabel metal2 s 37986 39200 38098 40000 6 io_out[6]
port 111 nsew signal bidirectional
rlabel metal3 s 0 15588 800 15828 6 io_out[7]
port 112 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 io_out[8]
port 113 nsew signal bidirectional
rlabel metal3 s 0 12188 800 12428 6 io_out[9]
port 114 nsew signal bidirectional
rlabel metal3 s 39200 6068 40000 6308 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 39200 4708 40000 4948 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 12870 39200 12982 40000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 25106 39200 25218 40000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 19310 39200 19422 40000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 14158 39200 14270 40000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 38630 39200 38742 40000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 39200 7428 40000 7668 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 39200 2668 40000 2908 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal2 s 634 39200 746 40000 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 33478 39200 33590 40000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 39200 19668 40000 19908 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 15446 39200 15558 40000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 16090 39200 16202 40000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_data_out[0]
port 147 nsew signal bidirectional
rlabel metal3 s 39200 9468 40000 9708 6 la1_data_out[10]
port 148 nsew signal bidirectional
rlabel metal2 s 18022 0 18134 800 6 la1_data_out[11]
port 149 nsew signal bidirectional
rlabel metal3 s 39200 36668 40000 36908 6 la1_data_out[12]
port 150 nsew signal bidirectional
rlabel metal2 s 3854 39200 3966 40000 6 la1_data_out[13]
port 151 nsew signal bidirectional
rlabel metal2 s 21242 39200 21354 40000 6 la1_data_out[14]
port 152 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal bidirectional
rlabel metal3 s 39200 13548 40000 13788 6 la1_data_out[16]
port 154 nsew signal bidirectional
rlabel metal3 s 39200 29188 40000 29428 6 la1_data_out[17]
port 155 nsew signal bidirectional
rlabel metal2 s 4498 39200 4610 40000 6 la1_data_out[18]
port 156 nsew signal bidirectional
rlabel metal3 s 39200 20348 40000 20588 6 la1_data_out[19]
port 157 nsew signal bidirectional
rlabel metal3 s 0 35988 800 36228 6 la1_data_out[1]
port 158 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 la1_data_out[20]
port 159 nsew signal bidirectional
rlabel metal3 s 39200 34628 40000 34868 6 la1_data_out[21]
port 160 nsew signal bidirectional
rlabel metal2 s 24462 39200 24574 40000 6 la1_data_out[22]
port 161 nsew signal bidirectional
rlabel metal2 s 9650 0 9762 800 6 la1_data_out[23]
port 162 nsew signal bidirectional
rlabel metal3 s 39200 14908 40000 15148 6 la1_data_out[24]
port 163 nsew signal bidirectional
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 164 nsew signal bidirectional
rlabel metal3 s 39200 4028 40000 4268 6 la1_data_out[26]
port 165 nsew signal bidirectional
rlabel metal3 s 0 38708 800 38948 6 la1_data_out[27]
port 166 nsew signal bidirectional
rlabel metal2 s 35410 0 35522 800 6 la1_data_out[28]
port 167 nsew signal bidirectional
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 168 nsew signal bidirectional
rlabel metal2 s 16734 0 16846 800 6 la1_data_out[2]
port 169 nsew signal bidirectional
rlabel metal3 s 39200 10148 40000 10388 6 la1_data_out[30]
port 170 nsew signal bidirectional
rlabel metal3 s 39200 38708 40000 38948 6 la1_data_out[31]
port 171 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[3]
port 172 nsew signal bidirectional
rlabel metal2 s 36698 0 36810 800 6 la1_data_out[4]
port 173 nsew signal bidirectional
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 174 nsew signal bidirectional
rlabel metal3 s 39200 16268 40000 16508 6 la1_data_out[6]
port 175 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal bidirectional
rlabel metal3 s 39200 29868 40000 30108 6 la1_data_out[8]
port 177 nsew signal bidirectional
rlabel metal2 s 37342 39200 37454 40000 6 la1_data_out[9]
port 178 nsew signal bidirectional
rlabel metal2 s 39274 0 39386 800 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 36054 39200 36166 40000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s 2566 39200 2678 40000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 17378 39200 17490 40000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 25750 39200 25862 40000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 16734 39200 16846 40000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 31546 39200 31658 40000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 39200 8108 40000 8348 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 39200 27828 40000 28068 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 6748 800 6988 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 39200 27148 40000 27388 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 22530 0 22642 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 27682 39200 27794 40000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 27038 39200 27150 40000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 5786 39200 5898 40000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 211 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 211 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 212 nsew ground input
rlabel metal3 s 39200 18988 40000 19228 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
