* NGSPICE file created from wrapped_cpr.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

.subckt wrapped_cpr active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12] la1_data_in[13] la1_data_in[14]
+ la1_data_in[15] la1_data_in[16] la1_data_in[17] la1_data_in[18] la1_data_in[19]
+ la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22] la1_data_in[23] la1_data_in[24]
+ la1_data_in[25] la1_data_in[26] la1_data_in[27] la1_data_in[28] la1_data_in[29]
+ la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3] la1_data_in[4] la1_data_in[5]
+ la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9] la1_data_out[0] la1_data_out[10]
+ la1_data_out[11] la1_data_out[12] la1_data_out[13] la1_data_out[14] la1_data_out[15]
+ la1_data_out[16] la1_data_out[17] la1_data_out[18] la1_data_out[19] la1_data_out[1]
+ la1_data_out[20] la1_data_out[21] la1_data_out[22] la1_data_out[23] la1_data_out[24]
+ la1_data_out[25] la1_data_out[26] la1_data_out[27] la1_data_out[28] la1_data_out[29]
+ la1_data_out[2] la1_data_out[30] la1_data_out[31] la1_data_out[3] la1_data_out[4]
+ la1_data_out[5] la1_data_out[6] la1_data_out[7] la1_data_out[8] la1_data_out[9]
+ la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12] la1_oenb[13] la1_oenb[14] la1_oenb[15]
+ la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19] la1_oenb[1] la1_oenb[20] la1_oenb[21]
+ la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25] la1_oenb[26] la1_oenb[27] la1_oenb[28]
+ la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31] la1_oenb[3] la1_oenb[4] la1_oenb[5]
+ la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9] vccd1 vssd1 wb_clk_i
X_2037_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2042_/A sky130_fd_sc_hd__buf_8
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2106_ _2549_/Q _2317_/A _2106_/C _2305_/A vssd1 vssd1 vccd1 vccd1 _2358_/B sky130_fd_sc_hd__and4_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1270_ _1270_/A _1514_/C _1438_/B vssd1 vssd1 vccd1 vccd1 _1278_/C sky130_fd_sc_hd__or3b_1
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1606_ _2493_/Q _1611_/A _1611_/C vssd1 vssd1 vccd1 vccd1 _1606_/X sky130_fd_sc_hd__and3_1
X_2724_ _2724_/A _2017_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1537_ _2494_/Q _2493_/Q _1611_/A _2487_/Q vssd1 vssd1 vccd1 vccd1 _1538_/D sky130_fd_sc_hd__and4_1
X_1468_ _1468_/A _1472_/D _1468_/C vssd1 vssd1 vccd1 vccd1 _1476_/A sky130_fd_sc_hd__and3_1
X_1399_ _1399_/A vssd1 vssd1 vccd1 vccd1 _2538_/D sky130_fd_sc_hd__clkinv_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2618__46 vssd1 vssd1 vccd1 vccd1 _2618__46/HI _2722_/A sky130_fd_sc_hd__conb_1
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2440_ _2544_/CLK _2440_/D _2163_/Y vssd1 vssd1 vccd1 vccd1 _2440_/Q sky130_fd_sc_hd__dfrtp_1
X_2632__60 vssd1 vssd1 vccd1 vccd1 _2632__60/HI _2740_/A sky130_fd_sc_hd__conb_1
X_1322_ _2549_/Q _2556_/Q _2555_/Q _2550_/Q vssd1 vssd1 vccd1 vccd1 _1323_/D sky130_fd_sc_hd__or4b_1
X_2371_ _2371_/A vssd1 vssd1 vccd1 vccd1 _2563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2569_ _2574_/CLK _2569_/D vssd1 vssd1 vccd1 vccd1 _2569_/Q sky130_fd_sc_hd__dfxtp_1
X_2707_ _2707_/A _1997_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1871_ _2436_/Q _1871_/B vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__or2_1
X_1940_ _1946_/A _1936_/C _2418_/Q vssd1 vssd1 vccd1 vccd1 _1940_/X sky130_fd_sc_hd__a21o_1
X_2423_ _2431_/CLK _2423_/D _2143_/Y vssd1 vssd1 vccd1 vccd1 _2423_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1305_ _1665_/C _1665_/D _1304_/Y vssd1 vssd1 vccd1 vccd1 _1847_/B sky130_fd_sc_hd__a21oi_2
X_2354_ _2560_/Q _2559_/Q _2354_/C vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__and3b_1
X_2285_ _2288_/A vssd1 vssd1 vccd1 vccd1 _2285_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2602__30 vssd1 vssd1 vccd1 vccd1 _2602__30/HI _2706_/A sky130_fd_sc_hd__conb_1
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2070_ _2072_/A vssd1 vssd1 vccd1 vccd1 _2070_/Y sky130_fd_sc_hd__inv_2
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1923_ _1933_/A _1923_/B vssd1 vssd1 vccd1 vccd1 _1923_/Y sky130_fd_sc_hd__nand2_1
X_1785_ _1785_/A _1789_/A vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__xor2_1
X_1854_ _1854_/A _1854_/B vssd1 vssd1 vccd1 vccd1 _1855_/A sky130_fd_sc_hd__and2_1
X_2406_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2573_/D sky130_fd_sc_hd__clkbuf_1
X_2199_ _2202_/A vssd1 vssd1 vccd1 vccd1 _2199_/Y sky130_fd_sc_hd__inv_2
X_2337_ _2344_/C vssd1 vssd1 vccd1 vccd1 _2337_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2575__3 vssd1 vssd1 vccd1 vccd1 _2575__3/HI _2679_/A sky130_fd_sc_hd__conb_1
X_2268_ _2270_/A vssd1 vssd1 vccd1 vccd1 _2268_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _2503_/Q _1570_/B vssd1 vssd1 vccd1 vccd1 _1577_/C sky130_fd_sc_hd__and2_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2053_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2053_/Y sky130_fd_sc_hd__inv_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _2122_/A vssd1 vssd1 vccd1 vccd1 _2410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2593__21 vssd1 vssd1 vccd1 vccd1 _2593__21/HI _2697_/A sky130_fd_sc_hd__conb_1
X_1906_ _1906_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__or2_1
X_1837_ _2439_/Q _1866_/A _2437_/Q _1872_/B vssd1 vssd1 vccd1 vccd1 _1847_/C sky130_fd_sc_hd__and4_1
X_1768_ _1765_/B _1767_/Y _2461_/Q _1676_/X vssd1 vssd1 vccd1 vccd1 _2461_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1699_ _1774_/B vssd1 vssd1 vccd1 vccd1 _1706_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1622_ _1634_/A _1625_/B _2490_/Q vssd1 vssd1 vccd1 vccd1 _1623_/C sky130_fd_sc_hd__a21oi_1
X_2740_ _2740_/A _2038_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1553_ _2507_/Q _1553_/B vssd1 vssd1 vccd1 vccd1 _1555_/C sky130_fd_sc_hd__nand2_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ _1484_/A _1658_/A vssd1 vssd1 vccd1 vccd1 _1484_/Y sky130_fd_sc_hd__nor2_1
X_2036_ input1/X vssd1 vssd1 vccd1 vccd1 _2061_/A sky130_fd_sc_hd__buf_2
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2105_ _2546_/Q _2545_/Q _2301_/C _2548_/Q vssd1 vssd1 vccd1 vccd1 _2305_/A sky130_fd_sc_hd__and4_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2723_ _2723_/A _2016_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_1536_ _2492_/Q vssd1 vssd1 vccd1 vccd1 _1611_/A sky130_fd_sc_hd__clkbuf_1
X_1605_ _1603_/Y _1608_/B _1595_/X _1657_/A vssd1 vssd1 vccd1 vccd1 _2495_/D sky130_fd_sc_hd__a211oi_1
XFILLER_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1467_ _1467_/A _1650_/A vssd1 vssd1 vccd1 vccd1 _1467_/Y sky130_fd_sc_hd__nand2_1
X_1398_ _1671_/A _1555_/B _1394_/Y _1397_/X vssd1 vssd1 vccd1 vccd1 _1399_/A sky130_fd_sc_hd__o31a_1
X_2019_ _2023_/A vssd1 vssd1 vccd1 vccd1 _2019_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2544_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_1321_ _2558_/Q _2557_/Q _2560_/Q _2559_/Q vssd1 vssd1 vccd1 vccd1 _1323_/C sky130_fd_sc_hd__or4_1
X_2370_ _2366_/X _2369_/Y _2563_/Q vssd1 vssd1 vccd1 vccd1 _2371_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2706_ _2706_/A _1996_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
X_2568_ _2568_/CLK _2568_/D vssd1 vssd1 vccd1 vccd1 _2568_/Q sky130_fd_sc_hd__dfxtp_1
X_1519_ _1519_/A _1519_/B _1519_/C _1519_/D vssd1 vssd1 vccd1 vccd1 _1519_/X sky130_fd_sc_hd__or4_1
X_2499_ _2522_/CLK _2499_/D _2237_/Y vssd1 vssd1 vccd1 vccd1 _2499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1870_ _1341_/X _1868_/Y _1869_/X _2437_/Q _1844_/X vssd1 vssd1 vccd1 vccd1 _2437_/D
+ sky130_fd_sc_hd__a32o_1
X_2422_ _2431_/CLK _2422_/D _2140_/Y vssd1 vssd1 vccd1 vccd1 _2422_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2353_ _2559_/Q _2354_/C _2352_/Y vssd1 vssd1 vccd1 vccd1 _2559_/D sky130_fd_sc_hd__o21a_1
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1304_ _2544_/Q _2543_/Q vssd1 vssd1 vccd1 vccd1 _1304_/Y sky130_fd_sc_hd__nand2_1
X_2284_ _2288_/A vssd1 vssd1 vccd1 vccd1 _2284_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1999_ _1999_/A vssd1 vssd1 vccd1 vccd1 _2004_/A sky130_fd_sc_hd__buf_8
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2669__97 vssd1 vssd1 vccd1 vccd1 _2669__97/HI _2777_/A sky130_fd_sc_hd__conb_1
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1922_ _1922_/A vssd1 vssd1 vccd1 vccd1 _2424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1784_ _1773_/A _1761_/X _1708_/A _1783_/X vssd1 vssd1 vccd1 vccd1 _2458_/D sky130_fd_sc_hd__a22o_1
X_1853_ _1307_/A _1847_/C _2440_/Q vssd1 vssd1 vccd1 vccd1 _1854_/B sky130_fd_sc_hd__a21o_1
X_2336_ _2336_/A _2336_/B _2555_/Q _2358_/B vssd1 vssd1 vccd1 vccd1 _2344_/C sky130_fd_sc_hd__and4_1
X_2405_ _2405_/A _2405_/B vssd1 vssd1 vccd1 vccd1 _2406_/A sky130_fd_sc_hd__and2_1
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2198_ _2202_/A vssd1 vssd1 vccd1 vccd1 _2198_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2267_ _2270_/A vssd1 vssd1 vccd1 vccd1 _2267_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2121_ _2121_/A _2121_/B vssd1 vssd1 vccd1 vccd1 _2122_/A sky130_fd_sc_hd__and2_1
X_2052_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2052_/Y sky130_fd_sc_hd__inv_2
X_1905_ _1905_/A vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1836_ _2436_/Q _2423_/Q _1908_/C _1836_/D vssd1 vssd1 vccd1 vccd1 _1872_/B sky130_fd_sc_hd__and4_1
X_1767_ _2461_/Q _1696_/A _1706_/A vssd1 vssd1 vccd1 vccd1 _1767_/Y sky130_fd_sc_hd__o21ai_1
X_1698_ _1848_/A _1698_/B vssd1 vssd1 vccd1 vccd1 _1774_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2319_ _2314_/A _2317_/A _2314_/B _2551_/Q vssd1 vssd1 vccd1 vccd1 _2319_/X sky130_fd_sc_hd__a31o_1
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2639__67 vssd1 vssd1 vccd1 vccd1 _2639__67/HI _2747_/A sky130_fd_sc_hd__conb_1
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1621_ _2491_/Q _1623_/B _1620_/Y vssd1 vssd1 vccd1 vccd1 _2491_/D sky130_fd_sc_hd__o21a_1
X_1552_ _1552_/A vssd1 vssd1 vccd1 vccd1 _2509_/D sky130_fd_sc_hd__clkbuf_1
X_2104_ _2547_/Q vssd1 vssd1 vccd1 vccd1 _2301_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1483_ _1483_/A vssd1 vssd1 vccd1 vccd1 _1483_/Y sky130_fd_sc_hd__inv_2
X_2035_ _2035_/A vssd1 vssd1 vccd1 vccd1 _2035_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2653__81 vssd1 vssd1 vccd1 vccd1 _2653__81/HI _2761_/A sky130_fd_sc_hd__conb_1
X_1819_ _1734_/A _1761_/A _2445_/Q vssd1 vssd1 vccd1 vccd1 _1820_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2722_ _2722_/A _2015_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1535_ _2491_/Q _2490_/Q _2489_/Q _2488_/Q vssd1 vssd1 vccd1 vccd1 _1563_/B sky130_fd_sc_hd__and4_1
X_1604_ _1633_/A _1604_/B vssd1 vssd1 vccd1 vccd1 _1608_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1466_ _1658_/A _1457_/C _1464_/Y _1465_/Y vssd1 vssd1 vccd1 vccd1 _2524_/D sky130_fd_sc_hd__o31ai_1
X_1397_ _1403_/A _1589_/A _1417_/A _1569_/A _1396_/Y vssd1 vssd1 vccd1 vccd1 _1397_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2018_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2023_/A sky130_fd_sc_hd__buf_4
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2609__37 vssd1 vssd1 vccd1 vccd1 _2609__37/HI _2713_/A sky130_fd_sc_hd__conb_1
XFILLER_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1320_ _2546_/Q _2545_/Q _2547_/Q _2548_/Q vssd1 vssd1 vccd1 vccd1 _1323_/B sky130_fd_sc_hd__or4b_2
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623__51 vssd1 vssd1 vccd1 vccd1 _2623__51/HI _2731_/A sky130_fd_sc_hd__conb_1
X_2705_ _2705_/A _1995_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
X_2567_ _2568_/CLK _2567_/D vssd1 vssd1 vccd1 vccd1 _2567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1449_ _1442_/B _1449_/B vssd1 vssd1 vccd1 vccd1 _1450_/A sky130_fd_sc_hd__and2b_1
X_1518_ _1669_/A _1669_/B _1669_/C _1518_/D vssd1 vssd1 vccd1 vccd1 _1519_/D sky130_fd_sc_hd__or4_1
X_2498_ _2522_/CLK _2498_/D _2236_/Y vssd1 vssd1 vccd1 vccd1 _2498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2421_ _2431_/CLK _2421_/D _2139_/Y vssd1 vssd1 vccd1 vccd1 _2421_/Q sky130_fd_sc_hd__dfrtp_1
X_2352_ _2352_/A _2352_/B vssd1 vssd1 vccd1 vccd1 _2352_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1303_ _1303_/A _1303_/B _1303_/C _1303_/D vssd1 vssd1 vccd1 vccd1 _1665_/D sky130_fd_sc_hd__nor4_2
X_2283_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2288_/A sky130_fd_sc_hd__buf_2
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1998_ _1998_/A vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__inv_2
X_2677__105 vssd1 vssd1 vccd1 vccd1 _2677__105/HI _2785_/A sky130_fd_sc_hd__conb_1
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1921_ _1921_/A _1921_/B vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__and2_1
X_1852_ _1852_/A vssd1 vssd1 vccd1 vccd1 _2441_/D sky130_fd_sc_hd__clkbuf_1
X_1783_ _1773_/A _1775_/X _1774_/C vssd1 vssd1 vccd1 vccd1 _1783_/X sky130_fd_sc_hd__o21ba_1
X_2335_ _2336_/A _2386_/A _2333_/B _2334_/Y vssd1 vssd1 vccd1 vccd1 _2554_/D sky130_fd_sc_hd__o31ai_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2404_ _2407_/A _2302_/A _2407_/D _2573_/Q vssd1 vssd1 vccd1 vccd1 _2405_/B sky130_fd_sc_hd__a31o_1
X_2266_ _2270_/A vssd1 vssd1 vccd1 vccd1 _2266_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2197_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2202_/A sky130_fd_sc_hd__buf_2
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2120_ _2407_/A _2112_/C _2399_/A _2407_/D _2410_/Q vssd1 vssd1 vccd1 vccd1 _2121_/B
+ sky130_fd_sc_hd__a41o_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2051_/Y sky130_fd_sc_hd__inv_2
X_1904_ _1341_/X _1901_/Y _1902_/X _1902_/A _1903_/X vssd1 vssd1 vccd1 vccd1 _2429_/D
+ sky130_fd_sc_hd__a32o_1
X_1835_ _1874_/B _1861_/A _1875_/B vssd1 vssd1 vccd1 vccd1 _1836_/D sky130_fd_sc_hd__and3_1
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1697_ _2474_/Q _2473_/Q _1716_/B vssd1 vssd1 vccd1 vccd1 _1704_/B sky130_fd_sc_hd__and3_1
X_1766_ _1734_/X _1763_/B _1765_/X _1755_/X _1765_/A vssd1 vssd1 vccd1 vccd1 _2462_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2318_ _2318_/A vssd1 vssd1 vccd1 vccd1 _2318_/Y sky130_fd_sc_hd__inv_2
X_2249_ _2252_/A vssd1 vssd1 vccd1 vccd1 _2249_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2584__12 vssd1 vssd1 vccd1 vccd1 _2584__12/HI _2688_/A sky130_fd_sc_hd__conb_1
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1620_ _1555_/B _1611_/C _1625_/A vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__o21ai_1
X_1551_ _1551_/A _1551_/B vssd1 vssd1 vccd1 vccd1 _1552_/A sky130_fd_sc_hd__and2_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1482_ _1451_/X _1480_/Y _1481_/X _1465_/B _1480_/A vssd1 vssd1 vccd1 vccd1 _2520_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2103_ _2552_/Q _2551_/Q vssd1 vssd1 vccd1 vccd1 _2106_/C sky130_fd_sc_hd__and2_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ _2035_/A vssd1 vssd1 vccd1 vccd1 _2034_/Y sky130_fd_sc_hd__inv_2
X_1818_ _1815_/B _1715_/A _1817_/X _1680_/X _2446_/Q vssd1 vssd1 vccd1 vccd1 _2446_/D
+ sky130_fd_sc_hd__a32o_1
X_1749_ _1749_/A vssd1 vssd1 vccd1 vccd1 _2467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2721_ _2721_/A _2014_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1534_ _2486_/Q _1638_/A _2484_/Q _2483_/Q vssd1 vssd1 vccd1 vccd1 _1562_/C sky130_fd_sc_hd__and4_1
X_1603_ _2495_/Q vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__inv_2
X_1465_ _1465_/A _1465_/B vssd1 vssd1 vccd1 vccd1 _1465_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1396_ _1671_/A vssd1 vssd1 vccd1 vccd1 _1396_/Y sky130_fd_sc_hd__inv_2
X_2017_ _2017_/A vssd1 vssd1 vccd1 vccd1 _2017_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2704_ _2704_/A _1994_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
X_2566_ _2566_/CLK _2566_/D vssd1 vssd1 vccd1 vccd1 _2566_/Q sky130_fd_sc_hd__dfxtp_1
X_2497_ _2506_/CLK _2497_/D _2233_/Y vssd1 vssd1 vccd1 vccd1 _2497_/Q sky130_fd_sc_hd__dfrtp_1
X_1448_ _1453_/A _1589_/A _1453_/B _1382_/A _2528_/Q vssd1 vssd1 vccd1 vccd1 _1449_/B
+ sky130_fd_sc_hd__a32o_1
X_1517_ _2536_/Q _1668_/A _2533_/Q _2535_/Q vssd1 vssd1 vccd1 vccd1 _1518_/D sky130_fd_sc_hd__or4bb_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1379_ _2540_/Q _1513_/A _1375_/B vssd1 vssd1 vccd1 vccd1 _1380_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2420_ _2431_/CLK _2420_/D _2138_/Y vssd1 vssd1 vccd1 vccd1 _2420_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2351_ _2109_/D _2350_/C _2386_/A vssd1 vssd1 vccd1 vccd1 _2352_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1302_ _2496_/Q _2495_/Q _2494_/Q _2493_/Q vssd1 vssd1 vccd1 vccd1 _1303_/D sky130_fd_sc_hd__or4_1
XFILLER_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2282_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2282_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ _1998_/A vssd1 vssd1 vccd1 vccd1 _1997_/Y sky130_fd_sc_hd__inv_2
X_2549_ _2574_/CLK _2549_/D vssd1 vssd1 vccd1 vccd1 _2549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1920_ _1925_/A _1885_/A _1908_/C _2424_/Q vssd1 vssd1 vccd1 vccd1 _1921_/B sky130_fd_sc_hd__a31o_1
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1851_ _1847_/X _1854_/A _2441_/Q vssd1 vssd1 vccd1 vccd1 _1852_/A sky130_fd_sc_hd__mux2_1
X_1782_ _1782_/A vssd1 vssd1 vccd1 vccd1 _2459_/D sky130_fd_sc_hd__clkbuf_1
X_2403_ _2403_/A _2403_/B vssd1 vssd1 vccd1 vccd1 _2405_/A sky130_fd_sc_hd__nand2_1
X_2196_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2196_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2334_ _2320_/A _2333_/X _2336_/A vssd1 vssd1 vccd1 vccd1 _2334_/Y sky130_fd_sc_hd__o21ai_1
X_2265_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2270_/A sky130_fd_sc_hd__buf_2
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2050_/Y sky130_fd_sc_hd__inv_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1834_ _2431_/Q _2430_/Q _2429_/Q _1906_/A vssd1 vssd1 vccd1 vccd1 _1875_/B sky130_fd_sc_hd__and4_1
X_1765_ _1765_/A _1765_/B vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__or2_1
X_1903_ _1903_/A vssd1 vssd1 vccd1 vccd1 _1903_/X sky130_fd_sc_hd__clkbuf_2
X_1696_ _1696_/A _1719_/C _1720_/C _1696_/D vssd1 vssd1 vccd1 vccd1 _1716_/B sky130_fd_sc_hd__and4_1
X_2179_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2184_/A sky130_fd_sc_hd__buf_2
X_2317_ _2317_/A _2551_/Q _2317_/C vssd1 vssd1 vccd1 vccd1 _2318_/A sky130_fd_sc_hd__and3_1
X_2248_ _2252_/A vssd1 vssd1 vccd1 vccd1 _2248_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1550_ _2508_/Q _2507_/Q _1577_/B _1553_/B _2509_/Q vssd1 vssd1 vccd1 vccd1 _1551_/B
+ sky130_fd_sc_hd__a41o_1
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2566_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1481_ _1483_/A _1455_/A _1455_/B _1480_/A vssd1 vssd1 vccd1 vccd1 _1481_/X sky130_fd_sc_hd__a31o_1
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2102_ _2550_/Q vssd1 vssd1 vccd1 vccd1 _2317_/A sky130_fd_sc_hd__clkbuf_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ _2035_/A vssd1 vssd1 vccd1 vccd1 _2033_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1817_ _2446_/Q _2445_/Q vssd1 vssd1 vccd1 vccd1 _1817_/X sky130_fd_sc_hd__or2_1
X_1748_ _1748_/A _1748_/B vssd1 vssd1 vccd1 vccd1 _1749_/A sky130_fd_sc_hd__and2_1
X_1679_ _1698_/B vssd1 vssd1 vccd1 vccd1 _1737_/B sky130_fd_sc_hd__buf_2
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2644__72 vssd1 vssd1 vccd1 vccd1 _2644__72/HI _2752_/A sky130_fd_sc_hd__conb_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1602_ _2496_/Q _1595_/X _1601_/Y vssd1 vssd1 vccd1 vccd1 _2496_/D sky130_fd_sc_hd__a21oi_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2720_ _2720_/A _2013_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
X_1533_ _2485_/Q vssd1 vssd1 vccd1 vccd1 _1638_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1464_ _1467_/A _1484_/A _1468_/C _1465_/A vssd1 vssd1 vccd1 vccd1 _1464_/Y sky130_fd_sc_hd__a31oi_1
X_1395_ _1468_/A vssd1 vssd1 vccd1 vccd1 _1589_/A sky130_fd_sc_hd__buf_2
X_2016_ _2017_/A vssd1 vssd1 vccd1 vccd1 _2016_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2565_ _2568_/CLK _2565_/D vssd1 vssd1 vccd1 vccd1 _2565_/Q sky130_fd_sc_hd__dfxtp_1
X_2703_ _2703_/A _1992_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_1516_ _2527_/Q _2522_/Q _2521_/Q _2528_/Q vssd1 vssd1 vccd1 vccd1 _1669_/C sky130_fd_sc_hd__or4b_1
X_2578__6 vssd1 vssd1 vccd1 vccd1 _2578__6/HI _2682_/A sky130_fd_sc_hd__conb_1
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2496_ _2506_/CLK _2496_/D _2232_/Y vssd1 vssd1 vccd1 vccd1 _2496_/Q sky130_fd_sc_hd__dfrtp_1
X_1447_ _1442_/A _1442_/B _1444_/X vssd1 vssd1 vccd1 vccd1 _2529_/D sky130_fd_sc_hd__o21a_1
X_1378_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1513_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2614__42 vssd1 vssd1 vccd1 vccd1 _2614__42/HI _2718_/A sky130_fd_sc_hd__conb_1
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2350_ _2558_/Q _2407_/C _2350_/C vssd1 vssd1 vccd1 vccd1 _2354_/C sky130_fd_sc_hd__and3_1
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1301_ _2488_/Q _2487_/Q _2486_/Q _2485_/Q vssd1 vssd1 vccd1 vccd1 _1303_/C sky130_fd_sc_hd__or4_1
X_2281_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2281_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _1998_/A vssd1 vssd1 vccd1 vccd1 _1996_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2548_ _2574_/CLK _2548_/D vssd1 vssd1 vccd1 vccd1 _2548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2479_ _2566_/CLK _2479_/D _2212_/Y vssd1 vssd1 vccd1 vccd1 _2479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2506_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1781_ _1781_/A _1781_/B vssd1 vssd1 vccd1 vccd1 _1782_/A sky130_fd_sc_hd__and2_1
X_1850_ _1878_/A _1850_/B vssd1 vssd1 vccd1 vccd1 _1854_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2333_ _2333_/A _2333_/B vssd1 vssd1 vccd1 vccd1 _2333_/X sky130_fd_sc_hd__and2_1
X_2402_ _2407_/A _2573_/Q _2119_/A _2393_/A vssd1 vssd1 vccd1 vccd1 _2403_/B sky130_fd_sc_hd__a31o_1
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2195_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2195_/Y sky130_fd_sc_hd__inv_2
X_2264_ _2264_/A vssd1 vssd1 vccd1 vccd1 _2264_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1979_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1979_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1902_ _1902_/A _1905_/A vssd1 vssd1 vccd1 vccd1 _1902_/X sky130_fd_sc_hd__or2_1
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1833_ _2428_/Q vssd1 vssd1 vccd1 vccd1 _1906_/A sky130_fd_sc_hd__clkbuf_1
X_1764_ _2463_/Q _1761_/X _1708_/A _1763_/Y vssd1 vssd1 vccd1 vccd1 _2463_/D sky130_fd_sc_hd__a22o_1
X_1695_ _2472_/Q _2471_/Q _2470_/Q _2469_/Q vssd1 vssd1 vccd1 vccd1 _1696_/D sky130_fd_sc_hd__and4_1
X_2316_ _2317_/A _2313_/Y _2315_/Y _2299_/X vssd1 vssd1 vccd1 vccd1 _2550_/D sky130_fd_sc_hd__o22a_1
X_2178_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2178_/Y sky130_fd_sc_hd__inv_2
X_2247_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2252_/A sky130_fd_sc_hd__buf_2
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1480_/A _1483_/A _1484_/A vssd1 vssd1 vccd1 vccd1 _1480_/Y sky130_fd_sc_hd__nand3_1
X_2032_ _2035_/A vssd1 vssd1 vccd1 vccd1 _2032_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2101_ _2561_/Q _2568_/Q _2382_/B _2374_/A vssd1 vssd1 vccd1 vccd1 _2110_/B sky130_fd_sc_hd__and4_1
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1678_ _2476_/Q vssd1 vssd1 vccd1 vccd1 _1678_/Y sky130_fd_sc_hd__inv_2
X_1816_ _2447_/Q _1755_/X _1715_/X _1815_/Y vssd1 vssd1 vccd1 vccd1 _2447_/D sky130_fd_sc_hd__a22o_1
X_1747_ _1734_/A _1751_/A _2467_/Q vssd1 vssd1 vccd1 vccd1 _1748_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1532_ _2482_/Q _2481_/Q _1654_/A _2479_/Q vssd1 vssd1 vccd1 vccd1 _1646_/B sky130_fd_sc_hd__and4_1
X_1601_ _2496_/Q _1595_/X _1503_/B vssd1 vssd1 vccd1 vccd1 _1601_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1463_ _1472_/D vssd1 vssd1 vccd1 vccd1 _1484_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1394_ _1403_/A _1417_/A vssd1 vssd1 vccd1 vccd1 _1394_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2015_ _2017_/A vssd1 vssd1 vccd1 vccd1 _2015_/Y sky130_fd_sc_hd__inv_2
X_2779_ _2779_/A _2083_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2702_ _2702_/A _1991_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
X_2564_ _2568_/CLK _2564_/D vssd1 vssd1 vccd1 vccd1 _2564_/Q sky130_fd_sc_hd__dfxtp_1
X_2495_ _2506_/CLK _2495_/D _2231_/Y vssd1 vssd1 vccd1 vccd1 _2495_/Q sky130_fd_sc_hd__dfrtp_1
X_1515_ _2526_/Q _2525_/Q _2524_/Q _2523_/Q vssd1 vssd1 vccd1 vccd1 _1669_/A sky130_fd_sc_hd__nand4_1
X_1377_ _1387_/A _2113_/A vssd1 vssd1 vccd1 vccd1 _1382_/A sky130_fd_sc_hd__or2_2
X_1446_ _1446_/A vssd1 vssd1 vccd1 vccd1 _2530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1300_ _2484_/Q _2482_/Q _2481_/Q _2483_/Q vssd1 vssd1 vccd1 vccd1 _1303_/B sky130_fd_sc_hd__or4bb_1
X_2280_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2280_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1995_ _1998_/A vssd1 vssd1 vccd1 vccd1 _1995_/Y sky130_fd_sc_hd__inv_2
X_2580__8 vssd1 vssd1 vccd1 vccd1 _2580__8/HI _2684_/A sky130_fd_sc_hd__conb_1
XFILLER_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2478_ _2544_/CLK _2478_/D _2211_/Y vssd1 vssd1 vccd1 vccd1 _2727_/A sky130_fd_sc_hd__dfrtp_1
X_2547_ _2574_/CLK _2547_/D vssd1 vssd1 vccd1 vccd1 _2547_/Q sky130_fd_sc_hd__dfxtp_1
X_1429_ _1423_/Y _1430_/A _1431_/S _1428_/X vssd1 vssd1 vccd1 vccd1 _2534_/D sky130_fd_sc_hd__a31o_1
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1780_ _1773_/A _1742_/A _1775_/X _2459_/Q vssd1 vssd1 vccd1 vccd1 _1781_/B sky130_fd_sc_hd__a31o_1
X_2332_ _2298_/X _2333_/B _2331_/X _2320_/X _2336_/B vssd1 vssd1 vccd1 vccd1 _2553_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2401_ _2401_/A vssd1 vssd1 vccd1 vccd1 _2572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2194_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2194_/Y sky130_fd_sc_hd__inv_2
X_2263_ _2264_/A vssd1 vssd1 vccd1 vccd1 _2263_/Y sky130_fd_sc_hd__inv_2
X_1978_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1978_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2665__93 vssd1 vssd1 vccd1 vccd1 _2665__93/HI _2773_/A sky130_fd_sc_hd__conb_1
X_1901_ _1902_/A _1905_/A vssd1 vssd1 vccd1 vccd1 _1901_/Y sky130_fd_sc_hd__nand2_1
X_1832_ _1857_/A _1936_/C _1858_/C _1923_/B vssd1 vssd1 vccd1 vccd1 _1908_/C sky130_fd_sc_hd__and4_1
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1694_ _2468_/Q _2467_/Q _2466_/Q _2465_/Q vssd1 vssd1 vccd1 vccd1 _1720_/C sky130_fd_sc_hd__and4_1
X_1763_ _2463_/Q _1763_/B vssd1 vssd1 vccd1 vccd1 _1763_/Y sky130_fd_sc_hd__xnor2_1
X_2315_ _1795_/X _2317_/C _2317_/A vssd1 vssd1 vccd1 vccd1 _2315_/Y sky130_fd_sc_hd__o21ai_1
X_2246_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2246_/Y sky130_fd_sc_hd__inv_2
X_2177_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2177_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2100_ _2562_/Q _2382_/A _2563_/Q vssd1 vssd1 vccd1 vccd1 _2374_/A sky130_fd_sc_hd__and3_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2590__18 vssd1 vssd1 vccd1 vccd1 _2590__18/HI _2694_/A sky130_fd_sc_hd__conb_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2031_ _2035_/A vssd1 vssd1 vccd1 vccd1 _2031_/Y sky130_fd_sc_hd__inv_2
X_1815_ _2447_/Q _1815_/B vssd1 vssd1 vccd1 vccd1 _1815_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1677_ _2726_/A _1743_/C _1676_/X vssd1 vssd1 vccd1 vccd1 _2477_/D sky130_fd_sc_hd__o21a_1
X_1746_ _1746_/A vssd1 vssd1 vccd1 vccd1 _2468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2229_ _2233_/A vssd1 vssd1 vccd1 vccd1 _2229_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2635__63 vssd1 vssd1 vccd1 vccd1 _2635__63/HI _2743_/A sky130_fd_sc_hd__conb_1
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1531_ _2480_/Q vssd1 vssd1 vccd1 vccd1 _1654_/A sky130_fd_sc_hd__clkbuf_1
X_1462_ _1457_/C _1459_/B _1459_/X _1457_/A vssd1 vssd1 vccd1 vccd1 _2525_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1600_ _1600_/A _1600_/B vssd1 vssd1 vccd1 vccd1 _2497_/D sky130_fd_sc_hd__nor2_1
X_1393_ _1413_/A _1419_/A _1393_/C _1393_/D vssd1 vssd1 vccd1 vccd1 _1417_/A sky130_fd_sc_hd__and4_1
XFILLER_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2014_ _2017_/A vssd1 vssd1 vccd1 vccd1 _2014_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2778_ _2778_/A _2082_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1729_ _1732_/A _1734_/A _1722_/D _2471_/Q vssd1 vssd1 vccd1 vccd1 _1730_/B sky130_fd_sc_hd__a31o_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2701_ _2701_/A _1990_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2563_ _2572_/CLK _2563_/D vssd1 vssd1 vccd1 vccd1 _2563_/Q sky130_fd_sc_hd__dfxtp_1
X_2494_ _2506_/CLK _2494_/D _2230_/Y vssd1 vssd1 vccd1 vccd1 _2494_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1445_ _1442_/X _1444_/X _1445_/S vssd1 vssd1 vccd1 vccd1 _1446_/A sky130_fd_sc_hd__mux2_1
X_1514_ _1671_/A _2537_/Q _1514_/C _1437_/X vssd1 vssd1 vccd1 vccd1 _1519_/C sky130_fd_sc_hd__or4b_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1376_ _2541_/Q _1380_/A _1372_/Y vssd1 vssd1 vccd1 vccd1 _2541_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2605__33 vssd1 vssd1 vccd1 vccd1 _2605__33/HI _2709_/A sky130_fd_sc_hd__conb_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _1998_/A vssd1 vssd1 vccd1 vccd1 _1994_/Y sky130_fd_sc_hd__inv_2
X_2477_ _2559_/CLK _2477_/D _2209_/Y vssd1 vssd1 vccd1 vccd1 _2726_/A sky130_fd_sc_hd__dfrtp_1
X_2546_ _2574_/CLK _2546_/D vssd1 vssd1 vccd1 vccd1 _2546_/Q sky130_fd_sc_hd__dfxtp_1
X_1428_ _1465_/B _1427_/Y _1668_/A vssd1 vssd1 vccd1 vccd1 _1428_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1359_ _2526_/Q _1457_/A _1465_/A _1467_/A vssd1 vssd1 vccd1 vccd1 _1362_/C sky130_fd_sc_hd__and4_1
XFILLER_50_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2400_ _2399_/X _2396_/Y _2407_/A vssd1 vssd1 vccd1 vccd1 _2401_/A sky130_fd_sc_hd__mux2_1
X_2331_ _2336_/B _2356_/A vssd1 vssd1 vccd1 vccd1 _2331_/X sky130_fd_sc_hd__or2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2262_ _2264_/A vssd1 vssd1 vccd1 vccd1 _2262_/Y sky130_fd_sc_hd__inv_2
X_2193_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2193_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2596__24 vssd1 vssd1 vccd1 vccd1 _2596__24/HI _2700_/A sky130_fd_sc_hd__conb_1
X_1977_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1977_/Y sky130_fd_sc_hd__inv_2
X_2529_ _2537_/CLK _2529_/D _2273_/Y vssd1 vssd1 vccd1 vccd1 _2529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1900_ _1307_/X _1897_/C _1899_/X _2430_/Q _1844_/X vssd1 vssd1 vccd1 vccd1 _2430_/D
+ sky130_fd_sc_hd__a32o_1
X_1831_ _2422_/Q _2421_/Q _2420_/Q vssd1 vssd1 vccd1 vccd1 _1923_/B sky130_fd_sc_hd__and3_1
X_1693_ _2464_/Q _2463_/Q _1765_/A _2461_/Q vssd1 vssd1 vccd1 vccd1 _1719_/C sky130_fd_sc_hd__and4_1
X_1762_ _1765_/A _1765_/B vssd1 vssd1 vccd1 vccd1 _1763_/B sky130_fd_sc_hd__nand2_1
X_2176_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__inv_2
X_2314_ _2314_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2317_/C sky130_fd_sc_hd__and2_1
X_2245_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2245_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2030_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2035_/A sky130_fd_sc_hd__clkbuf_8
X_2673__101 vssd1 vssd1 vccd1 vccd1 _2673__101/HI _2781_/A sky130_fd_sc_hd__conb_1
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1814_ _1715_/A _1812_/Y _1813_/X _1680_/X _2448_/Q vssd1 vssd1 vccd1 vccd1 _2448_/D
+ sky130_fd_sc_hd__a32o_1
X_1745_ _1742_/X _1748_/A _2468_/Q vssd1 vssd1 vccd1 vccd1 _1746_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1676_ _1761_/A vssd1 vssd1 vccd1 vccd1 _1676_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2159_ _2159_/A vssd1 vssd1 vccd1 vccd1 _2159_/Y sky130_fd_sc_hd__inv_2
X_2228_ _2228_/A vssd1 vssd1 vccd1 vccd1 _2233_/A sky130_fd_sc_hd__buf_2
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2650__78 vssd1 vssd1 vccd1 vccd1 _2650__78/HI _2758_/A sky130_fd_sc_hd__conb_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1530_ _2502_/Q _2501_/Q _1591_/S _2495_/Q vssd1 vssd1 vccd1 vccd1 _1539_/B sky130_fd_sc_hd__and4_1
XFILLER_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1461_ _1461_/A vssd1 vssd1 vccd1 vccd1 _2526_/D sky130_fd_sc_hd__clkbuf_1
X_1392_ _1668_/B _1435_/A _1435_/B _1434_/A vssd1 vssd1 vccd1 vccd1 _1393_/D sky130_fd_sc_hd__and4_1
X_2013_ _2017_/A vssd1 vssd1 vccd1 vccd1 _2013_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1728_ _1728_/A vssd1 vssd1 vccd1 vccd1 _2472_/D sky130_fd_sc_hd__clkbuf_1
X_2777_ _2777_/A _2081_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ _1659_/A vssd1 vssd1 vccd1 vccd1 _1659_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2526_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2700_ _2700_/A _1989_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2562_ _2568_/CLK _2562_/D vssd1 vssd1 vccd1 vccd1 _2562_/Q sky130_fd_sc_hd__dfxtp_1
X_2493_ _2506_/CLK _2493_/D _2229_/Y vssd1 vssd1 vccd1 vccd1 _2493_/Q sky130_fd_sc_hd__dfrtp_1
X_1375_ _2540_/Q _1375_/B vssd1 vssd1 vccd1 vccd1 _1380_/A sky130_fd_sc_hd__and2_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1444_ _1444_/A _1444_/B vssd1 vssd1 vccd1 vccd1 _1444_/X sky130_fd_sc_hd__or2_1
X_1513_ _1513_/A vssd1 vssd1 vccd1 vccd1 _1643_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2620__48 vssd1 vssd1 vccd1 vccd1 _2620__48/HI _2724_/A sky130_fd_sc_hd__conb_1
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1998_/A sky130_fd_sc_hd__buf_6
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2545_ _2574_/CLK _2545_/D vssd1 vssd1 vccd1 vccd1 _2545_/Q sky130_fd_sc_hd__dfxtp_1
X_2476_ _2476_/CLK _2476_/D _2208_/Y vssd1 vssd1 vccd1 vccd1 _2476_/Q sky130_fd_sc_hd__dfrtp_1
X_1358_ _2523_/Q vssd1 vssd1 vccd1 vccd1 _1467_/A sky130_fd_sc_hd__clkbuf_1
X_1427_ _1430_/A _1393_/D _1658_/A vssd1 vssd1 vccd1 vccd1 _1427_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1289_ _1289_/A _1289_/B _1289_/C _1289_/D vssd1 vssd1 vccd1 vccd1 _1289_/X sky130_fd_sc_hd__or4_4
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2192_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2192_/Y sky130_fd_sc_hd__inv_2
X_2330_ _2336_/B _2356_/A vssd1 vssd1 vccd1 vccd1 _2333_/B sky130_fd_sc_hd__nand2_1
X_2261_ _2264_/A vssd1 vssd1 vccd1 vccd1 _2261_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1976_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1976_/Y sky130_fd_sc_hd__inv_2
X_2528_ _2537_/CLK _2528_/D _2272_/Y vssd1 vssd1 vccd1 vccd1 _2528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2459_ _2560_/CLK _2459_/D _2187_/Y vssd1 vssd1 vccd1 vccd1 _2459_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1761_ _1761_/A vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__clkbuf_2
X_1830_ _2419_/Q _2418_/Q vssd1 vssd1 vccd1 vccd1 _1858_/C sky130_fd_sc_hd__and2_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1692_ _2462_/Q vssd1 vssd1 vccd1 vccd1 _1765_/A sky130_fd_sc_hd__clkbuf_1
X_2313_ _2313_/A _2386_/A vssd1 vssd1 vccd1 vccd1 _2313_/Y sky130_fd_sc_hd__nor2_1
X_2175_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2175_/Y sky130_fd_sc_hd__inv_2
X_2244_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2244_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2522_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_2656__84 vssd1 vssd1 vccd1 vccd1 _2656__84/HI _2764_/A sky130_fd_sc_hd__conb_1
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _1959_/A vssd1 vssd1 vccd1 vccd1 _2412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1813_ _2447_/Q _2446_/Q _2445_/Q _2448_/Q vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__a31o_1
X_1744_ _1795_/A _1742_/B _1777_/A vssd1 vssd1 vccd1 vccd1 _1748_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1675_ _1698_/B vssd1 vssd1 vccd1 vccd1 _1761_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2158_ _2159_/A vssd1 vssd1 vccd1 vccd1 _2158_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2089_ _2090_/A vssd1 vssd1 vccd1 vccd1 _2089_/Y sky130_fd_sc_hd__inv_2
X_2227_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2227_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1460_ _1457_/X _1459_/X _2526_/Q vssd1 vssd1 vccd1 vccd1 _1461_/A sky130_fd_sc_hd__mux2_1
X_1391_ _1445_/S _1442_/A _1438_/B vssd1 vssd1 vccd1 vccd1 _1435_/B sky130_fd_sc_hd__and3_1
X_2012_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2017_/A sky130_fd_sc_hd__buf_6
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2626__54 vssd1 vssd1 vccd1 vccd1 _2626__54/HI _2734_/A sky130_fd_sc_hd__conb_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2776_ _2776_/A _2080_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_1727_ _1722_/X _1730_/A _2472_/Q vssd1 vssd1 vccd1 vccd1 _1728_/A sky130_fd_sc_hd__mux2_1
X_1658_ _1658_/A _1658_/B vssd1 vssd1 vccd1 vccd1 _1658_/Y sky130_fd_sc_hd__nor2_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1589_ _1589_/A _1589_/B _1595_/A vssd1 vssd1 vccd1 vccd1 _1589_/X sky130_fd_sc_hd__and3_1
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2561_ _2572_/CLK _2561_/D vssd1 vssd1 vccd1 vccd1 _2561_/Q sky130_fd_sc_hd__dfxtp_1
X_2492_ _2506_/CLK _2492_/D _2227_/Y vssd1 vssd1 vccd1 vccd1 _2492_/Q sky130_fd_sc_hd__dfrtp_1
X_1512_ _1512_/A vssd1 vssd1 vccd1 vccd1 _2511_/D sky130_fd_sc_hd__clkbuf_1
X_1374_ _1374_/A vssd1 vssd1 vccd1 vccd1 _2542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1443_ _1442_/A _1425_/C _1416_/A vssd1 vssd1 vccd1 vccd1 _1444_/B sky130_fd_sc_hd__a21oi_1
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2759_ _2759_/A _2059_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1992_ _1992_/A vssd1 vssd1 vccd1 vccd1 _1992_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2475_ _2476_/CLK _2475_/D _2207_/Y vssd1 vssd1 vccd1 vccd1 _2475_/Q sky130_fd_sc_hd__dfrtp_1
X_2544_ _2544_/CLK _2544_/D _2290_/Y vssd1 vssd1 vccd1 vccd1 _2544_/Q sky130_fd_sc_hd__dfrtp_1
X_1288_ _1288_/A _1288_/B _1288_/C _1288_/D vssd1 vssd1 vccd1 vccd1 _1289_/D sky130_fd_sc_hd__or4_1
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1357_ _2524_/Q vssd1 vssd1 vccd1 vccd1 _1465_/A sky130_fd_sc_hd__clkbuf_1
X_1426_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1465_/B sky130_fd_sc_hd__buf_2
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2191_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2196_/A sky130_fd_sc_hd__buf_2
X_2260_ _2264_/A vssd1 vssd1 vccd1 vccd1 _2260_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1980_/A sky130_fd_sc_hd__buf_8
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2458_ _2560_/CLK _2458_/D _2186_/Y vssd1 vssd1 vccd1 vccd1 _2458_/Q sky130_fd_sc_hd__dfrtp_1
X_2527_ _2537_/CLK _2527_/D _2270_/Y vssd1 vssd1 vccd1 vccd1 _2527_/Q sky130_fd_sc_hd__dfrtp_1
X_1409_ _1409_/A _1409_/B _1409_/C _1669_/B vssd1 vssd1 vccd1 vccd1 _1409_/X sky130_fd_sc_hd__or4_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2389_ _2399_/A _2393_/B _2115_/A vssd1 vssd1 vccd1 vccd1 _2391_/A sky130_fd_sc_hd__a21o_1
X_2587__15 vssd1 vssd1 vccd1 vccd1 _2587__15/HI _2691_/A sky130_fd_sc_hd__conb_1
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1760_ _1734_/X _1757_/Y _1759_/X _1755_/X _2464_/Q vssd1 vssd1 vccd1 vccd1 _2464_/D
+ sky130_fd_sc_hd__a32o_1
X_1691_ _1800_/A _1758_/C vssd1 vssd1 vccd1 vccd1 _1696_/A sky130_fd_sc_hd__and2_1
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2312_ _2313_/A _2302_/X _2311_/X _2299_/X _2314_/A vssd1 vssd1 vccd1 vccd1 _2549_/D
+ sky130_fd_sc_hd__a32o_1
X_2174_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2174_/Y sky130_fd_sc_hd__inv_2
X_2243_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2243_/Y sky130_fd_sc_hd__inv_2
X_2671__99 vssd1 vssd1 vccd1 vccd1 _2671__99/HI _2779_/A sky130_fd_sc_hd__conb_1
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1889_ _1889_/A vssd1 vssd1 vccd1 vccd1 _2433_/D sky130_fd_sc_hd__clkbuf_1
X_1958_ _1885_/A _1903_/A _1958_/S vssd1 vssd1 vccd1 vccd1 _1959_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1812_ _1812_/A vssd1 vssd1 vccd1 vccd1 _1812_/Y sky130_fd_sc_hd__inv_2
X_1743_ _1886_/A _1743_/B _1743_/C vssd1 vssd1 vccd1 vccd1 _1777_/A sky130_fd_sc_hd__and3_1
X_1674_ _1710_/A _1710_/B _1743_/B _1743_/C vssd1 vssd1 vccd1 vccd1 _1698_/B sky130_fd_sc_hd__o211ai_4
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2226_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2226_/Y sky130_fd_sc_hd__inv_2
X_2088_ _2090_/A vssd1 vssd1 vccd1 vccd1 _2088_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2157_ _2159_/A vssd1 vssd1 vccd1 vccd1 _2157_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ _2529_/Q vssd1 vssd1 vccd1 vccd1 _1442_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2011_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2011_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2641__69 vssd1 vssd1 vccd1 vccd1 _2641__69/HI _2749_/A sky130_fd_sc_hd__conb_1
X_2775_ _2775_/A _2078_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_1726_ _1737_/B _1726_/B vssd1 vssd1 vccd1 vccd1 _1730_/A sky130_fd_sc_hd__or2_1
X_1657_ _1657_/A _1657_/B _1657_/C vssd1 vssd1 vccd1 vccd1 _2480_/D sky130_fd_sc_hd__nor3_1
X_1588_ _1588_/A vssd1 vssd1 vccd1 vccd1 _2501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _2209_/A vssd1 vssd1 vccd1 vccd1 _2209_/Y sky130_fd_sc_hd__inv_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2560_ _2560_/CLK _2560_/D vssd1 vssd1 vccd1 vccd1 _2560_/Q sky130_fd_sc_hd__dfxtp_1
X_2491_ _2491_/CLK _2491_/D _2226_/Y vssd1 vssd1 vccd1 vccd1 _2491_/Q sky130_fd_sc_hd__dfrtp_1
X_1442_ _1442_/A _1442_/B vssd1 vssd1 vccd1 vccd1 _1442_/X sky130_fd_sc_hd__and2_1
X_1511_ _1451_/X _1459_/A _1511_/S vssd1 vssd1 vccd1 vccd1 _1512_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1373_ _1372_/B _1372_/Y _2542_/Q vssd1 vssd1 vccd1 vccd1 _1374_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2758_ _2758_/A _2058_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
X_1709_ _1704_/B _1708_/Y _2474_/Q _1676_/X vssd1 vssd1 vccd1 vccd1 _2474_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2689_ _2689_/A _1976_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_64_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2611__39 vssd1 vssd1 vccd1 vccd1 _2611__39/HI _2715_/A sky130_fd_sc_hd__conb_1
X_1991_ _1992_/A vssd1 vssd1 vccd1 vccd1 _1991_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2474_ _2476_/CLK _2474_/D _2206_/Y vssd1 vssd1 vccd1 vccd1 _2474_/Q sky130_fd_sc_hd__dfrtp_1
X_2543_ _2559_/CLK _2543_/D _2289_/Y vssd1 vssd1 vccd1 vccd1 _2543_/Q sky130_fd_sc_hd__dfrtp_1
X_1425_ _1468_/A _1425_/B _1425_/C vssd1 vssd1 vccd1 vccd1 _1431_/S sky130_fd_sc_hd__and3_1
X_1287_ _2450_/Q _2449_/Q _2447_/Q _2448_/Q vssd1 vssd1 vccd1 vccd1 _1288_/D sky130_fd_sc_hd__or4b_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1356_ _2525_/Q vssd1 vssd1 vccd1 vccd1 _1457_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ _2190_/A vssd1 vssd1 vccd1 vccd1 _2190_/Y sky130_fd_sc_hd__inv_2
X_1974_ input1/X vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__buf_2
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2457_ _2560_/CLK _2457_/D _2184_/Y vssd1 vssd1 vccd1 vccd1 _2457_/Q sky130_fd_sc_hd__dfrtp_1
X_2388_ _2388_/A vssd1 vssd1 vccd1 vccd1 _2568_/D sky130_fd_sc_hd__clkbuf_1
X_2526_ _2526_/CLK _2526_/D _2269_/Y vssd1 vssd1 vccd1 vccd1 _2526_/Q sky130_fd_sc_hd__dfrtp_1
X_1408_ _2516_/Q _2515_/Q _2520_/Q _2519_/Q vssd1 vssd1 vccd1 vccd1 _1669_/B sky130_fd_sc_hd__or4bb_1
X_1339_ _1339_/A _1339_/B _1339_/C _1339_/D vssd1 vssd1 vccd1 vccd1 _1710_/B sky130_fd_sc_hd__nor4_4
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1690_ _2460_/Q _1690_/B _1690_/C vssd1 vssd1 vccd1 vccd1 _1758_/C sky130_fd_sc_hd__and3_1
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2311_ _2314_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__or2_1
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2242_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2242_/Y sky130_fd_sc_hd__inv_2
X_2173_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2178_/A sky130_fd_sc_hd__buf_2
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ _1821_/X _1333_/D _1956_/Y _1956_/A _1824_/X vssd1 vssd1 vccd1 vccd1 _2413_/D
+ sky130_fd_sc_hd__a32o_1
X_1888_ _1885_/X _1891_/A _2433_/Q vssd1 vssd1 vccd1 vccd1 _1889_/A sky130_fd_sc_hd__mux2_1
X_2509_ _2566_/CLK _2509_/D _2249_/Y vssd1 vssd1 vccd1 vccd1 _2509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2647__75 vssd1 vssd1 vccd1 vccd1 _2647__75/HI _2755_/A sky130_fd_sc_hd__conb_1
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1811_ _1715_/A _1803_/B _1810_/X _1680_/X _2449_/Q vssd1 vssd1 vccd1 vccd1 _2449_/D
+ sky130_fd_sc_hd__a32o_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1742_ _1742_/A _1742_/B vssd1 vssd1 vccd1 vccd1 _1742_/X sky130_fd_sc_hd__and2_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1673_ _1669_/X _1672_/X _1259_/A vssd1 vssd1 vccd1 vccd1 _1743_/C sky130_fd_sc_hd__o21ai_4
X_2225_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2225_/Y sky130_fd_sc_hd__inv_2
X_2156_ _2159_/A vssd1 vssd1 vccd1 vccd1 _2156_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2087_ _2090_/A vssd1 vssd1 vccd1 vccd1 _2087_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2010_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1725_ _1732_/B _1723_/Y _2333_/A vssd1 vssd1 vccd1 vccd1 _1726_/B sky130_fd_sc_hd__o21a_1
X_2774_ _2774_/A _2077_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1656_ _1659_/A _1634_/A _1654_/A vssd1 vssd1 vccd1 vccd1 _1657_/C sky130_fd_sc_hd__a21oi_1
X_1587_ _1643_/A _1587_/B _1587_/C vssd1 vssd1 vccd1 vccd1 _1588_/A sky130_fd_sc_hd__and3_1
X_2208_ _2209_/A vssd1 vssd1 vccd1 vccd1 _2208_/Y sky130_fd_sc_hd__inv_2
X_2139_ _2140_/A vssd1 vssd1 vccd1 vccd1 _2139_/Y sky130_fd_sc_hd__inv_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2617__45 vssd1 vssd1 vccd1 vccd1 _2617__45/HI _2721_/A sky130_fd_sc_hd__conb_1
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2490_ _2491_/CLK _2490_/D _2225_/Y vssd1 vssd1 vccd1 vccd1 _2490_/Q sky130_fd_sc_hd__dfrtp_1
X_1510_ _1501_/A _1509_/X _1505_/Y _1465_/B _1509_/A vssd1 vssd1 vccd1 vccd1 _2512_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1441_ _1435_/A _1439_/X _1436_/X vssd1 vssd1 vccd1 vccd1 _2531_/D sky130_fd_sc_hd__o21a_1
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1372_ _1569_/A _1372_/B vssd1 vssd1 vccd1 vccd1 _1372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2688_ _2688_/A _1973_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
X_1708_ _1708_/A _1708_/B vssd1 vssd1 vccd1 vccd1 _1708_/Y sky130_fd_sc_hd__nand2_1
X_2757_ _2757_/A _2057_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_58_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1639_ _1639_/A _1639_/B _1639_/C vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__nand3_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1990_ _1992_/A vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2542_ _2568_/CLK _2542_/D _2288_/Y vssd1 vssd1 vccd1 vccd1 _2542_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2476_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_2473_ _2559_/CLK _2473_/D _2205_/Y vssd1 vssd1 vccd1 vccd1 _2473_/Q sky130_fd_sc_hd__dfrtp_1
X_1424_ _1438_/B _1434_/A vssd1 vssd1 vccd1 vccd1 _1425_/C sky130_fd_sc_hd__and2_1
X_1355_ _2518_/Q _1670_/D _1498_/S _1493_/A vssd1 vssd1 vccd1 vccd1 _1455_/B sky130_fd_sc_hd__and4_1
X_1286_ _2454_/Q _2453_/Q _2452_/Q _2451_/Q vssd1 vssd1 vccd1 vccd1 _1288_/C sky130_fd_sc_hd__or4_1
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1973_ _1973_/A vssd1 vssd1 vccd1 vccd1 _1973_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2525_ _2526_/CLK _2525_/D _2268_/Y vssd1 vssd1 vccd1 vccd1 _2525_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2456_ _2464_/CLK _2456_/D _2183_/Y vssd1 vssd1 vccd1 vccd1 _2456_/Q sky130_fd_sc_hd__dfrtp_1
X_1338_ _1338_/A _1338_/B _1874_/B _1861_/A vssd1 vssd1 vccd1 vccd1 _1339_/D sky130_fd_sc_hd__or4bb_1
X_2387_ _2386_/Y _2384_/B _2568_/Q vssd1 vssd1 vccd1 vccd1 _2388_/A sky130_fd_sc_hd__mux2_1
X_1407_ _2522_/Q _2517_/Q _2518_/Q _1472_/A vssd1 vssd1 vccd1 vccd1 _1409_/C sky130_fd_sc_hd__or4bb_1
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1269_ _2528_/Q _2527_/Q vssd1 vssd1 vccd1 vccd1 _1438_/B sky130_fd_sc_hd__and2_1
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2172_ _2234_/A vssd1 vssd1 vccd1 vccd1 _2197_/A sky130_fd_sc_hd__clkbuf_2
X_2310_ _2314_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2313_/A sky130_fd_sc_hd__nand2_1
X_2241_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2246_/A sky130_fd_sc_hd__buf_2
XFILLER_53_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1887_ _1911_/B _1885_/B _1795_/A vssd1 vssd1 vccd1 vccd1 _1891_/A sky130_fd_sc_hd__o21ai_1
X_1956_ _1956_/A _1958_/S vssd1 vssd1 vccd1 vccd1 _1956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2592__20 vssd1 vssd1 vccd1 vccd1 _2592__20/HI _2696_/A sky130_fd_sc_hd__conb_1
X_2508_ _2566_/CLK _2508_/D _2248_/Y vssd1 vssd1 vccd1 vccd1 _2508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2439_ _2439_/CLK _2439_/D _2162_/Y vssd1 vssd1 vccd1 vccd1 _2439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ _2449_/Q _1812_/A vssd1 vssd1 vccd1 vccd1 _1810_/X sky130_fd_sc_hd__or2_1
X_1741_ _2467_/Q _1751_/A vssd1 vssd1 vccd1 vccd1 _1742_/B sky130_fd_sc_hd__and2_1
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1672_ _1672_/A _1672_/B _1672_/C _1672_/D vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__or4_1
X_2155_ _2159_/A vssd1 vssd1 vccd1 vccd1 _2155_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2224_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2224_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2086_ _2090_/A vssd1 vssd1 vccd1 vccd1 _2086_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _1939_/A vssd1 vssd1 vccd1 vccd1 _1939_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2773_ _2773_/A _2076_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_1724_ _2113_/A vssd1 vssd1 vccd1 vccd1 _2333_/A sky130_fd_sc_hd__buf_2
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ _1625_/A _1653_/X _1657_/B _2481_/Q vssd1 vssd1 vccd1 vccd1 _2481_/D sky130_fd_sc_hd__o2bb2a_1
X_1586_ _1591_/S _1589_/B _1595_/A _2501_/Q vssd1 vssd1 vccd1 vccd1 _1587_/C sky130_fd_sc_hd__a31o_1
X_2069_ _2072_/A vssd1 vssd1 vccd1 vccd1 _2069_/Y sky130_fd_sc_hd__inv_2
X_2207_ _2209_/A vssd1 vssd1 vccd1 vccd1 _2207_/Y sky130_fd_sc_hd__inv_2
X_2138_ _2140_/A vssd1 vssd1 vccd1 vccd1 _2138_/Y sky130_fd_sc_hd__inv_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1440_ _1668_/B _1436_/X _1437_/X _1439_/X vssd1 vssd1 vccd1 vccd1 _2532_/D sky130_fd_sc_hd__a22o_1
X_1371_ _1584_/A vssd1 vssd1 vccd1 vccd1 _1569_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2756_ _2756_/A _2056_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_1707_ _2473_/Q _1716_/B _2474_/Q vssd1 vssd1 vccd1 vccd1 _1708_/B sky130_fd_sc_hd__a21o_1
X_2687_ _2687_/A _1972_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
X_1638_ _1638_/A vssd1 vssd1 vccd1 vccd1 _1638_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1569_ _1569_/A vssd1 vssd1 vccd1 vccd1 _1637_/A sky130_fd_sc_hd__clkbuf_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2472_ _2559_/CLK _2472_/D _2202_/Y vssd1 vssd1 vccd1 vccd1 _2472_/Q sky130_fd_sc_hd__dfrtp_1
X_2541_ _2568_/CLK _2541_/D _2287_/Y vssd1 vssd1 vccd1 vccd1 _2541_/Q sky130_fd_sc_hd__dfrtp_1
X_1285_ _2462_/Q _2461_/Q _2460_/Q _2459_/Q vssd1 vssd1 vccd1 vccd1 _1288_/B sky130_fd_sc_hd__or4_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1423_ _1668_/A vssd1 vssd1 vccd1 vccd1 _1423_/Y sky130_fd_sc_hd__inv_2
X_1354_ _2517_/Q vssd1 vssd1 vccd1 vccd1 _1670_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2739_ _2739_/A _2035_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2668__96 vssd1 vssd1 vccd1 vccd1 _2668__96/HI _2776_/A sky130_fd_sc_hd__conb_1
XFILLER_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1972_ _1973_/A vssd1 vssd1 vccd1 vccd1 _1972_/Y sky130_fd_sc_hd__inv_2
X_2455_ _2464_/CLK _2455_/D _2182_/Y vssd1 vssd1 vccd1 vccd1 _2455_/Q sky130_fd_sc_hd__dfrtp_1
X_2524_ _2526_/CLK _2524_/D _2267_/Y vssd1 vssd1 vccd1 vccd1 _2524_/Q sky130_fd_sc_hd__dfrtp_1
X_1337_ _2435_/Q _2434_/Q _2433_/Q _2432_/Q vssd1 vssd1 vccd1 vccd1 _1861_/A sky130_fd_sc_hd__and4_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2386_ _2386_/A _2386_/B vssd1 vssd1 vccd1 vccd1 _2386_/Y sky130_fd_sc_hd__nor2_1
X_1406_ _1668_/B _2531_/Q _2530_/Q _2529_/Q vssd1 vssd1 vccd1 vccd1 _1409_/B sky130_fd_sc_hd__nand4_1
X_1268_ _2518_/Q _2517_/Q vssd1 vssd1 vccd1 vccd1 _1514_/C sky130_fd_sc_hd__nand2_1
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2171_ _2171_/A vssd1 vssd1 vccd1 vccd1 _2171_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2240_ _2240_/A vssd1 vssd1 vccd1 vccd1 _2240_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1886_ _1886_/A vssd1 vssd1 vccd1 vccd1 _1911_/B sky130_fd_sc_hd__clkbuf_2
X_1955_ _1821_/X _1953_/Y _1954_/X _1953_/A _1824_/X vssd1 vssd1 vccd1 vccd1 _2414_/D
+ sky130_fd_sc_hd__a32o_1
X_2438_ _2544_/CLK _2438_/D _2161_/Y vssd1 vssd1 vccd1 vccd1 _2438_/Q sky130_fd_sc_hd__dfrtp_1
X_2507_ _2566_/CLK _2507_/D _2246_/Y vssd1 vssd1 vccd1 vccd1 _2507_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2369_ _2393_/A _2372_/C _2403_/A vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2638__66 vssd1 vssd1 vccd1 vccd1 _2638__66/HI _2746_/A sky130_fd_sc_hd__conb_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1740_ _2466_/Q _1754_/A _1740_/C vssd1 vssd1 vccd1 vccd1 _1751_/A sky130_fd_sc_hd__and3_1
XFILLER_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1671_ _1671_/A _2537_/Q _2530_/Q _2529_/Q vssd1 vssd1 vccd1 vccd1 _1672_/D sky130_fd_sc_hd__or4bb_1
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2085_ _2085_/A vssd1 vssd1 vccd1 vccd1 _2090_/A sky130_fd_sc_hd__buf_6
X_2154_ _2166_/A vssd1 vssd1 vccd1 vccd1 _2159_/A sky130_fd_sc_hd__buf_2
XFILLER_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2223_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2223_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2652__80 vssd1 vssd1 vccd1 vccd1 _2652__80/HI _2760_/A sky130_fd_sc_hd__conb_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1869_ _2437_/Q _1872_/B vssd1 vssd1 vccd1 vccd1 _1869_/X sky130_fd_sc_hd__or2_1
X_1938_ _1341_/X _1934_/B _1937_/X _2419_/Q _1903_/X vssd1 vssd1 vccd1 vccd1 _2419_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2772_ _2772_/A _2075_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
X_1723_ _2471_/Q _1732_/A vssd1 vssd1 vccd1 vccd1 _1723_/Y sky130_fd_sc_hd__nand2_1
X_1654_ _1654_/A _1659_/A _1654_/C vssd1 vssd1 vccd1 vccd1 _1657_/B sky130_fd_sc_hd__and3_1
X_2206_ _2209_/A vssd1 vssd1 vccd1 vccd1 _2206_/Y sky130_fd_sc_hd__inv_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _1582_/Y _1587_/B _1580_/X _1657_/A vssd1 vssd1 vccd1 vccd1 _2502_/D sky130_fd_sc_hd__a211oi_1
X_2137_ _2140_/A vssd1 vssd1 vccd1 vccd1 _2137_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2068_ _2072_/A vssd1 vssd1 vccd1 vccd1 _2068_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2608__36 vssd1 vssd1 vccd1 vccd1 _2608__36/HI _2712_/A sky130_fd_sc_hd__conb_1
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1370_ _2114_/A _2113_/A vssd1 vssd1 vccd1 vccd1 _1584_/A sky130_fd_sc_hd__nor2_2
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2622__50 vssd1 vssd1 vccd1 vccd1 _2622__50/HI _2730_/A sky130_fd_sc_hd__conb_1
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1706_ _1706_/A vssd1 vssd1 vccd1 vccd1 _1708_/A sky130_fd_sc_hd__clkbuf_2
X_1637_ _1637_/A _1637_/B _1636_/X vssd1 vssd1 vccd1 vccd1 _2486_/D sky130_fd_sc_hd__nor3b_1
X_2755_ _2755_/A _2054_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
X_2686_ _2686_/A _1971_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1568_ _2507_/Q _1572_/B _1554_/X vssd1 vssd1 vccd1 vccd1 _2507_/D sky130_fd_sc_hd__o21a_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1499_/A vssd1 vssd1 vccd1 vccd1 _2516_/D sky130_fd_sc_hd__clkbuf_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2471_ _2559_/CLK _2471_/D _2201_/Y vssd1 vssd1 vccd1 vccd1 _2471_/Q sky130_fd_sc_hd__dfrtp_1
X_2540_ _2572_/CLK _2540_/D _2286_/Y vssd1 vssd1 vccd1 vccd1 _2540_/Q sky130_fd_sc_hd__dfrtp_1
X_1422_ _1422_/A vssd1 vssd1 vccd1 vccd1 _2535_/D sky130_fd_sc_hd__inv_2
X_1284_ _2458_/Q _2457_/Q _2456_/Q _2455_/Q vssd1 vssd1 vccd1 vccd1 _1288_/A sky130_fd_sc_hd__or4_1
X_1353_ _2514_/Q _2513_/Q _1509_/A _1511_/S vssd1 vssd1 vccd1 vccd1 _1455_/A sky130_fd_sc_hd__and4_1
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2599__27 vssd1 vssd1 vccd1 vccd1 _2599__27/HI _2703_/A sky130_fd_sc_hd__conb_1
X_2738_ _2738_/A _2034_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2676__104 vssd1 vssd1 vccd1 vccd1 _2676__104/HI _2784_/A sky130_fd_sc_hd__conb_1
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ _1973_/A vssd1 vssd1 vccd1 vccd1 _1971_/Y sky130_fd_sc_hd__inv_2
X_2454_ _2464_/CLK _2454_/D _2181_/Y vssd1 vssd1 vccd1 vccd1 _2454_/Q sky130_fd_sc_hd__dfrtp_1
X_2385_ _2566_/Q _2378_/X _2386_/B _2384_/X vssd1 vssd1 vccd1 vccd1 _2567_/D sky130_fd_sc_hd__a31o_1
X_2523_ _2526_/CLK _2523_/D _2266_/Y vssd1 vssd1 vccd1 vccd1 _2523_/Q sky130_fd_sc_hd__dfrtp_1
X_1405_ _1419_/A _1420_/B _1413_/A vssd1 vssd1 vccd1 vccd1 _1417_/B sky130_fd_sc_hd__a21oi_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
X_1336_ _2427_/Q _2426_/Q _2425_/Q _2424_/Q vssd1 vssd1 vccd1 vccd1 _1874_/B sky130_fd_sc_hd__and4_1
XFILLER_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1267_ _2524_/Q _2523_/Q vssd1 vssd1 vccd1 vccd1 _1270_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2170_ _2171_/A vssd1 vssd1 vccd1 vccd1 _2170_/Y sky130_fd_sc_hd__inv_2
X_1954_ _1956_/A _1958_/S _1953_/A vssd1 vssd1 vccd1 vccd1 _1954_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1885_ _1885_/A _1885_/B vssd1 vssd1 vccd1 vccd1 _1885_/X sky130_fd_sc_hd__and2_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2437_ _2439_/CLK _2437_/D _2159_/Y vssd1 vssd1 vccd1 vccd1 _2437_/Q sky130_fd_sc_hd__dfrtp_1
X_2368_ _2381_/A _2563_/Q _2374_/C vssd1 vssd1 vccd1 vccd1 _2372_/C sky130_fd_sc_hd__and3_1
X_2506_ _2506_/CLK _2506_/D _2245_/Y vssd1 vssd1 vccd1 vccd1 _2506_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2299_ _2320_/A vssd1 vssd1 vccd1 vccd1 _2299_/X sky130_fd_sc_hd__clkbuf_2
X_1319_ _2562_/Q _2561_/Q _2564_/Q _2563_/Q vssd1 vssd1 vccd1 vccd1 _1323_/A sky130_fd_sc_hd__or4_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2583__11 vssd1 vssd1 vccd1 vccd1 _2583__11/HI _2687_/A sky130_fd_sc_hd__conb_1
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1670_ _2536_/Q _2535_/Q _2518_/Q _1670_/D vssd1 vssd1 vccd1 vccd1 _1672_/C sky130_fd_sc_hd__nand4b_1
X_2222_ _2228_/A vssd1 vssd1 vccd1 vccd1 _2227_/A sky130_fd_sc_hd__buf_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_2153_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2153_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ _2084_/A vssd1 vssd1 vccd1 vccd1 _2084_/Y sky130_fd_sc_hd__inv_2
X_1937_ _2419_/Q _1939_/A vssd1 vssd1 vccd1 vccd1 _1937_/X sky130_fd_sc_hd__or2_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1799_ _1734_/X _1794_/Y _1798_/X _1755_/X _1798_/A vssd1 vssd1 vccd1 vccd1 _2453_/D
+ sky130_fd_sc_hd__a32o_1
X_1868_ _1868_/A vssd1 vssd1 vccd1 vccd1 _1868_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2771_ _2771_/A _2074_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
X_1722_ _2471_/Q _1732_/A _1742_/A _1722_/D vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__and4_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1653_ _2481_/Q _1654_/A _1659_/A _1555_/B vssd1 vssd1 vccd1 vccd1 _1653_/X sky130_fd_sc_hd__a31o_1
X_1584_ _1584_/A vssd1 vssd1 vccd1 vccd1 _1657_/A sky130_fd_sc_hd__buf_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2209_/A vssd1 vssd1 vccd1 vccd1 _2205_/Y sky130_fd_sc_hd__inv_2
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2067_ _2085_/A vssd1 vssd1 vccd1 vccd1 _2072_/A sky130_fd_sc_hd__buf_8
X_2136_ _2140_/A vssd1 vssd1 vccd1 vccd1 _2136_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1705_ _2475_/Q _1703_/X _1700_/Y _1704_/X vssd1 vssd1 vccd1 vccd1 _2475_/D sky130_fd_sc_hd__a22o_1
X_2754_ _2754_/A _2053_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1636_ _1638_/A _1639_/A _1633_/A _1639_/C _2486_/Q vssd1 vssd1 vccd1 vccd1 _1636_/X
+ sky130_fd_sc_hd__a41o_1
X_2685_ _2685_/A _1970_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
X_1567_ _1567_/A _1580_/A _1593_/C vssd1 vssd1 vccd1 vccd1 _1572_/B sky130_fd_sc_hd__and3_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2119_ _2119_/A vssd1 vssd1 vccd1 vccd1 _2407_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1497_/B _1497_/Y _1498_/S vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__mux2_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2470_ _2559_/CLK _2470_/D _2200_/Y vssd1 vssd1 vccd1 vccd1 _2470_/Q sky130_fd_sc_hd__dfrtp_1
X_1421_ _1419_/A _1419_/Y _1421_/S vssd1 vssd1 vccd1 vccd1 _1422_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1283_ _2470_/Q _2469_/Q _2468_/Q _2467_/Q vssd1 vssd1 vccd1 vccd1 _1289_/C sky130_fd_sc_hd__or4_1
X_1352_ _2511_/Q vssd1 vssd1 vccd1 vccd1 _1511_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_2737_ _2737_/A _2033_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
X_1619_ _2490_/Q _1654_/C _1625_/B vssd1 vssd1 vccd1 vccd1 _1623_/B sky130_fd_sc_hd__and3_1
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1970_ _1973_/A vssd1 vssd1 vccd1 vccd1 _1970_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2522_ _2522_/CLK _2522_/D _2264_/Y vssd1 vssd1 vccd1 vccd1 _2522_/Q sky130_fd_sc_hd__dfrtp_2
X_2453_ _2464_/CLK _2453_/D _2180_/Y vssd1 vssd1 vccd1 vccd1 _2453_/Q sky130_fd_sc_hd__dfrtp_1
X_1335_ _2421_/Q _2420_/Q _2418_/Q _2419_/Q vssd1 vssd1 vccd1 vccd1 _1338_/B sky130_fd_sc_hd__or4b_1
X_2384_ _2567_/Q _2384_/B vssd1 vssd1 vccd1 vccd1 _2384_/X sky130_fd_sc_hd__and2_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1404_ _1403_/A _1402_/X _1403_/X _1501_/A vssd1 vssd1 vccd1 vccd1 _2537_/D sky130_fd_sc_hd__a22o_1
X_2659__87 vssd1 vssd1 vccd1 vccd1 _2659__87/HI _2767_/A sky130_fd_sc_hd__conb_1
Xinput2 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
X_1266_ _1445_/S _2529_/Q vssd1 vssd1 vccd1 vccd1 _1519_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2559_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1884_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1885_/A sky130_fd_sc_hd__clkbuf_2
X_1953_ _1953_/A _1956_/A _1958_/S vssd1 vssd1 vccd1 vccd1 _1953_/Y sky130_fd_sc_hd__nand3_1
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2505_ _2566_/CLK _2505_/D _2244_/Y vssd1 vssd1 vccd1 vccd1 _2505_/Q sky130_fd_sc_hd__dfrtp_1
X_2576__4 vssd1 vssd1 vccd1 vccd1 _2576__4/HI _2680_/A sky130_fd_sc_hd__conb_1
XFILLER_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2436_ _2439_/CLK _2436_/D _2158_/Y vssd1 vssd1 vccd1 vccd1 _2436_/Q sky130_fd_sc_hd__dfrtp_1
X_2367_ _2367_/A vssd1 vssd1 vccd1 vccd1 _2393_/A sky130_fd_sc_hd__clkbuf_2
X_2298_ _2302_/A vssd1 vssd1 vccd1 vccd1 _2298_/X sky130_fd_sc_hd__clkbuf_2
X_1318_ _1318_/A _1318_/B _1318_/C _1318_/D vssd1 vssd1 vccd1 vccd1 _2113_/B sky130_fd_sc_hd__nor4_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2152_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2152_/Y sky130_fd_sc_hd__inv_2
X_2221_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2221_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2083_ _2084_/A vssd1 vssd1 vccd1 vccd1 _2083_/Y sky130_fd_sc_hd__inv_2
X_2629__57 vssd1 vssd1 vccd1 vccd1 _2629__57/HI _2737_/A sky130_fd_sc_hd__conb_1
X_1936_ _2418_/Q _1946_/A _1936_/C vssd1 vssd1 vccd1 vccd1 _1939_/A sky130_fd_sc_hd__and3_1
X_1867_ _1844_/X _1866_/A _1863_/Y _1866_/X vssd1 vssd1 vccd1 vccd1 _2438_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1798_ _1798_/A _1800_/A vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__or2_1
X_2419_ _2431_/CLK _2419_/D _2137_/Y vssd1 vssd1 vccd1 vccd1 _2419_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2643__71 vssd1 vssd1 vccd1 vccd1 _2643__71/HI _2751_/A sky130_fd_sc_hd__conb_1
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2770_ _2770_/A _2072_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_1721_ _1732_/B vssd1 vssd1 vccd1 vccd1 _1722_/D sky130_fd_sc_hd__inv_2
XFILLER_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ _2479_/Q vssd1 vssd1 vccd1 vccd1 _1659_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1583_ _2501_/Q _1591_/S _1589_/B _1593_/C vssd1 vssd1 vccd1 vccd1 _1587_/B sky130_fd_sc_hd__nand4_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _2290_/A vssd1 vssd1 vccd1 vccd1 _2140_/A sky130_fd_sc_hd__buf_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2228_/A vssd1 vssd1 vccd1 vccd1 _2209_/A sky130_fd_sc_hd__buf_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2066_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2066_/Y sky130_fd_sc_hd__inv_2
X_1919_ _1919_/A vssd1 vssd1 vccd1 vccd1 _2425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1704_ _2475_/Q _1704_/B vssd1 vssd1 vccd1 vccd1 _1704_/X sky130_fd_sc_hd__or2_1
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2684_ _2684_/A _1969_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
X_2753_ _2753_/A _2052_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_1635_ _2487_/Q _1637_/B _1634_/Y _1503_/B vssd1 vssd1 vccd1 vccd1 _2487_/D sky130_fd_sc_hd__o211a_1
X_1566_ _1595_/A vssd1 vssd1 vccd1 vccd1 _1593_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1569_/A _1497_/B vssd1 vssd1 vccd1 vccd1 _1497_/Y sky130_fd_sc_hd__nor2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__buf_8
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2118_ _2407_/C vssd1 vssd1 vccd1 vccd1 _2399_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2613__41 vssd1 vssd1 vccd1 vccd1 _2613__41/HI _2717_/A sky130_fd_sc_hd__conb_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1351_ _2512_/Q vssd1 vssd1 vccd1 vccd1 _1509_/A sky130_fd_sc_hd__clkbuf_1
X_1420_ _1589_/A _1420_/B vssd1 vssd1 vccd1 vccd1 _1421_/S sky130_fd_sc_hd__nand2_1
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1282_ _2466_/Q _2465_/Q _2464_/Q _2463_/Q vssd1 vssd1 vccd1 vccd1 _1289_/B sky130_fd_sc_hd__or4_1
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2736_ _2736_/A _2032_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
X_1618_ _2489_/Q _2488_/Q _1634_/B vssd1 vssd1 vccd1 vccd1 _1625_/B sky130_fd_sc_hd__and3_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1549_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1577_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ _2526_/CLK _2521_/D _2263_/Y vssd1 vssd1 vccd1 vccd1 _2521_/Q sky130_fd_sc_hd__dfrtp_1
X_2452_ _2464_/CLK _2452_/D _2178_/Y vssd1 vssd1 vccd1 vccd1 _2452_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1334_ _2417_/Q _2416_/Q _2415_/Q _2414_/Q vssd1 vssd1 vccd1 vccd1 _1338_/A sky130_fd_sc_hd__or4_1
X_2383_ _2124_/B _2386_/B _2115_/A vssd1 vssd1 vccd1 vccd1 _2384_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1265_ _2530_/Q vssd1 vssd1 vccd1 vccd1 _1445_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_1403_ _1403_/A _1417_/A vssd1 vssd1 vccd1 vccd1 _1403_/X sky130_fd_sc_hd__xor2_1
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2719_ _2719_/A _2011_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1883_ _1883_/A vssd1 vssd1 vccd1 vccd1 _2434_/D sky130_fd_sc_hd__clkbuf_1
X_1952_ _1821_/X _1947_/B _1951_/X _2415_/Q _1903_/X vssd1 vssd1 vccd1 vccd1 _2415_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2435_ _2559_/CLK _2435_/D _2157_/Y vssd1 vssd1 vccd1 vccd1 _2435_/Q sky130_fd_sc_hd__dfrtp_1
X_2504_ _2566_/CLK _2504_/D _2243_/Y vssd1 vssd1 vccd1 vccd1 _2504_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1317_ _2552_/Q _2551_/Q _2336_/A _2553_/Q vssd1 vssd1 vccd1 vccd1 _1318_/D sky130_fd_sc_hd__nand4_1
X_2297_ _2301_/A _2301_/B vssd1 vssd1 vccd1 vccd1 _2297_/Y sky130_fd_sc_hd__nand2_1
X_2366_ _2381_/A _2399_/A _2382_/D vssd1 vssd1 vccd1 vccd1 _2366_/X sky130_fd_sc_hd__and3_1
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2151_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2151_/Y sky130_fd_sc_hd__inv_2
X_2082_ _2084_/A vssd1 vssd1 vccd1 vccd1 _2082_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2220_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2220_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1797_ _1787_/B _1796_/X _2454_/Q _1676_/X vssd1 vssd1 vccd1 vccd1 _2454_/D sky130_fd_sc_hd__a2bb2o_1
X_1935_ _2420_/Q _1934_/Y _1930_/X vssd1 vssd1 vccd1 vccd1 _2420_/D sky130_fd_sc_hd__o21a_1
X_1866_ _1866_/A _1868_/A vssd1 vssd1 vccd1 vccd1 _1866_/X sky130_fd_sc_hd__or2_1
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2418_ _2491_/CLK _2418_/D _2136_/Y vssd1 vssd1 vccd1 vccd1 _2418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2349_ _2349_/A _2349_/B vssd1 vssd1 vccd1 vccd1 _2558_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1720_ _2469_/Q _1740_/C _1720_/C vssd1 vssd1 vccd1 vccd1 _1732_/B sky130_fd_sc_hd__nand3_2
X_1651_ _1651_/A vssd1 vssd1 vccd1 vccd1 _2482_/D sky130_fd_sc_hd__clkbuf_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _2502_/Q vssd1 vssd1 vccd1 vccd1 _1582_/Y sky130_fd_sc_hd__inv_2
X_2065_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2065_/Y sky130_fd_sc_hd__inv_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _2134_/A vssd1 vssd1 vccd1 vccd1 _2134_/Y sky130_fd_sc_hd__inv_2
X_2203_ _2234_/A vssd1 vssd1 vccd1 vccd1 _2228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1918_ _1916_/X _1921_/A _2425_/Q vssd1 vssd1 vccd1 vccd1 _1919_/A sky130_fd_sc_hd__mux2_1
X_1849_ _2440_/Q _1847_/C _1928_/A vssd1 vssd1 vccd1 vccd1 _1850_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1703_ _1761_/A vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__clkbuf_2
X_1634_ _1634_/A _1634_/B vssd1 vssd1 vccd1 vccd1 _1634_/Y sky130_fd_sc_hd__nand2_1
X_2683_ _2683_/A _1967_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
X_2752_ _2752_/A _2051_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_1565_ _1416_/A _1658_/B _1521_/Y _1564_/X vssd1 vssd1 vccd1 vccd1 _1595_/A sky130_fd_sc_hd__o211a_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1496_/A vssd1 vssd1 vccd1 vccd1 _2517_/D sky130_fd_sc_hd__inv_2
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2117_ _2572_/Q vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2048_ _2048_/A vssd1 vssd1 vccd1 vccd1 _2048_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1281_ _2476_/Q _2475_/Q _1281_/C _1815_/B vssd1 vssd1 vccd1 vccd1 _1289_/A sky130_fd_sc_hd__or4_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_1350_ _1668_/B _1435_/A _1445_/S _2529_/Q vssd1 vssd1 vccd1 vccd1 _1425_/B sky130_fd_sc_hd__and4_1
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1617_ _1617_/A vssd1 vssd1 vccd1 vccd1 _2492_/D sky130_fd_sc_hd__clkbuf_1
X_2735_ _2735_/A _2031_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1548_ _1474_/X _1544_/C _1547_/X vssd1 vssd1 vccd1 vccd1 _1551_/A sky130_fd_sc_hd__o21ai_1
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1479_ _1451_/X _1473_/Y _1478_/X _1402_/X _1472_/A vssd1 vssd1 vccd1 vccd1 _2521_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2451_ _2464_/CLK _2451_/D _2177_/Y vssd1 vssd1 vccd1 vccd1 _2451_/Q sky130_fd_sc_hd__dfrtp_1
X_1402_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1402_/X sky130_fd_sc_hd__clkbuf_2
X_2520_ _2522_/CLK _2520_/D _2262_/Y vssd1 vssd1 vccd1 vccd1 _2520_/Q sky130_fd_sc_hd__dfrtp_1
X_1333_ _2443_/Q _2442_/Q _1333_/C _1333_/D vssd1 vssd1 vccd1 vccd1 _1339_/C sky130_fd_sc_hd__or4_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2382_ _2382_/A _2382_/B _2382_/C _2382_/D vssd1 vssd1 vccd1 vccd1 _2386_/B sky130_fd_sc_hd__nand4_2
X_1264_ _1672_/A _1672_/B vssd1 vssd1 vccd1 vccd1 _1519_/A sky130_fd_sc_hd__or2_1
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2718_ _2718_/A _2010_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2664__92 vssd1 vssd1 vccd1 vccd1 _2664__92/HI _2772_/A sky130_fd_sc_hd__conb_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1882_ _1881_/X _1878_/Y _2434_/Q vssd1 vssd1 vccd1 vccd1 _1883_/A sky130_fd_sc_hd__mux2_1
X_1951_ _1953_/A _1956_/A _1958_/S _2415_/Q vssd1 vssd1 vccd1 vccd1 _1951_/X sky130_fd_sc_hd__a31o_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2434_ _2476_/CLK _2434_/D _2156_/Y vssd1 vssd1 vccd1 vccd1 _2434_/Q sky130_fd_sc_hd__dfrtp_1
X_2365_ _2365_/A _2365_/B vssd1 vssd1 vccd1 vccd1 _2562_/D sky130_fd_sc_hd__nor2_1
X_2503_ _2506_/CLK _2503_/D _2242_/Y vssd1 vssd1 vccd1 vccd1 _2503_/Q sky130_fd_sc_hd__dfrtp_1
X_1316_ _2554_/Q vssd1 vssd1 vccd1 vccd1 _2336_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2296_ _2546_/Q vssd1 vssd1 vccd1 vccd1 _2301_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2150_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2150_/Y sky130_fd_sc_hd__inv_2
X_2081_ _2084_/A vssd1 vssd1 vccd1 vccd1 _2081_/Y sky130_fd_sc_hd__inv_2
X_1934_ _1947_/A _1934_/B vssd1 vssd1 vccd1 vccd1 _1934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1796_ _1793_/Y _1794_/Y _1737_/B _1795_/X vssd1 vssd1 vccd1 vccd1 _1796_/X sky130_fd_sc_hd__a211o_1
X_1865_ _1824_/X _1856_/Y _1863_/Y _1864_/X vssd1 vssd1 vccd1 vccd1 _2439_/D sky130_fd_sc_hd__o31a_1
X_2417_ _2491_/CLK _2417_/D _2134_/Y vssd1 vssd1 vccd1 vccd1 _2417_/Q sky130_fd_sc_hd__dfrtp_1
X_2348_ _1878_/A _2350_/C _2352_/A _2558_/Q vssd1 vssd1 vccd1 vccd1 _2349_/B sky130_fd_sc_hd__o211a_1
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2279_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2279_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2634__62 vssd1 vssd1 vccd1 vccd1 _2634__62/HI _2742_/A sky130_fd_sc_hd__conb_1
X_1650_ _1650_/A _1650_/B _1650_/C vssd1 vssd1 vccd1 vccd1 _1651_/A sky130_fd_sc_hd__and3_1
X_1581_ _2503_/Q _1580_/X _1574_/Y vssd1 vssd1 vccd1 vccd1 _2503_/D sky130_fd_sc_hd__o21a_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2202_/A vssd1 vssd1 vccd1 vccd1 _2202_/Y sky130_fd_sc_hd__inv_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2133_ _2134_/A vssd1 vssd1 vccd1 vccd1 _2133_/Y sky130_fd_sc_hd__inv_2
X_2064_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2064_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1917_ _1911_/B _1916_/B _1795_/A vssd1 vssd1 vccd1 vccd1 _1921_/A sky130_fd_sc_hd__o21ai_1
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1779_ _1779_/A vssd1 vssd1 vccd1 vccd1 _2460_/D sky130_fd_sc_hd__clkbuf_1
X_1848_ _1848_/A vssd1 vssd1 vccd1 vccd1 _1878_/A sky130_fd_sc_hd__buf_2
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2751_ _2751_/A _2050_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1702_ _1678_/Y _1680_/X _1700_/Y _1701_/X vssd1 vssd1 vccd1 vccd1 _2476_/D sky130_fd_sc_hd__o31a_1
X_1633_ _1633_/A _1633_/B _1639_/C vssd1 vssd1 vccd1 vccd1 _1637_/B sky130_fd_sc_hd__and3_1
X_1564_ _2495_/Q _1564_/B _1611_/C vssd1 vssd1 vccd1 vccd1 _1564_/X sky130_fd_sc_hd__and3_1
X_2682_ _2682_/A _1966_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1670_/D _1490_/Y _1495_/S vssd1 vssd1 vccd1 vccd1 _1496_/A sky130_fd_sc_hd__mux2_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ _2048_/A vssd1 vssd1 vccd1 vccd1 _2047_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2116_ _2302_/A _2126_/B _2320_/A vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__a21o_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2604__32 vssd1 vssd1 vccd1 vccd1 _2604__32/HI _2708_/A sky130_fd_sc_hd__conb_1
X_1280_ _2446_/Q _2445_/Q vssd1 vssd1 vccd1 vccd1 _1815_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2734_ _2734_/A _2029_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1547_ _1612_/A vssd1 vssd1 vccd1 vccd1 _1547_/X sky130_fd_sc_hd__clkbuf_2
X_1616_ _1643_/A _1616_/B _1616_/C vssd1 vssd1 vccd1 vccd1 _1617_/A sky130_fd_sc_hd__and3_1
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1478_ _1480_/A _1483_/A _1484_/A _1472_/A vssd1 vssd1 vccd1 vccd1 _1478_/X sky130_fd_sc_hd__a31o_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2450_ _2464_/CLK _2450_/D _2176_/Y vssd1 vssd1 vccd1 vccd1 _2450_/Q sky130_fd_sc_hd__dfrtp_1
X_2381_ _2381_/A _2563_/Q vssd1 vssd1 vccd1 vccd1 _2382_/C sky130_fd_sc_hd__and2_1
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1401_ _1444_/A vssd1 vssd1 vccd1 vccd1 _1459_/A sky130_fd_sc_hd__clkbuf_2
X_1332_ _2413_/Q _2412_/Q vssd1 vssd1 vccd1 vccd1 _1333_/D sky130_fd_sc_hd__or2_1
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1263_ _2542_/Q _2541_/Q _2512_/Q _2511_/Q vssd1 vssd1 vccd1 vccd1 _1672_/B sky130_fd_sc_hd__or4_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2717_ _2717_/A _2009_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_2595__23 vssd1 vssd1 vccd1 vccd1 _2595__23/HI _2699_/A sky130_fd_sc_hd__conb_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1950_ _2412_/Q vssd1 vssd1 vccd1 vccd1 _1958_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1881_ _2433_/Q _1916_/A _1885_/B vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__and3_1
X_2502_ _2522_/CLK _2502_/D _2240_/Y vssd1 vssd1 vccd1 vccd1 _2502_/Q sky130_fd_sc_hd__dfrtp_1
X_2433_ _2476_/CLK _2433_/D _2155_/Y vssd1 vssd1 vccd1 vccd1 _2433_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2364_ _2302_/X _2382_/D _2381_/A vssd1 vssd1 vccd1 vccd1 _2365_/B sky130_fd_sc_hd__a21oi_1
X_1315_ _2574_/Q _2573_/Q _2411_/Q _2410_/Q vssd1 vssd1 vccd1 vccd1 _1318_/C sky130_fd_sc_hd__or4_1
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2295_ _2546_/Q _2545_/Q vssd1 vssd1 vccd1 vccd1 _2295_/X sky130_fd_sc_hd__or2_1
XFILLER_2_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ _2084_/A vssd1 vssd1 vccd1 vccd1 _2080_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1933_ _1933_/A vssd1 vssd1 vccd1 vccd1 _1934_/B sky130_fd_sc_hd__inv_2
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2464_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_1864_ _1866_/A _1307_/A _1868_/A _2439_/Q vssd1 vssd1 vccd1 vccd1 _1864_/X sky130_fd_sc_hd__a31o_1
X_1795_ _1795_/A vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__clkbuf_2
X_2416_ _2491_/CLK _2416_/D _2133_/Y vssd1 vssd1 vccd1 vccd1 _2416_/Q sky130_fd_sc_hd__dfrtp_1
X_2347_ _2372_/B _2350_/C _2558_/Q vssd1 vssd1 vccd1 vccd1 _2349_/A sky130_fd_sc_hd__a21oi_1
X_2672__100 vssd1 vssd1 vccd1 vccd1 _2672__100/HI _2780_/A sky130_fd_sc_hd__conb_1
X_2278_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2278_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1580_ _1580_/A _1593_/C vssd1 vssd1 vccd1 vccd1 _1580_/X sky130_fd_sc_hd__and2_1
X_2201_ _2202_/A vssd1 vssd1 vccd1 vccd1 _2201_/Y sky130_fd_sc_hd__inv_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _2134_/A vssd1 vssd1 vccd1 vccd1 _2132_/Y sky130_fd_sc_hd__inv_2
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2063_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2063_/Y sky130_fd_sc_hd__inv_2
X_1916_ _1916_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__and2_1
X_1847_ _2440_/Q _1847_/B _1847_/C vssd1 vssd1 vccd1 vccd1 _1847_/X sky130_fd_sc_hd__and3_1
X_1778_ _1774_/X _1781_/A _2460_/Q vssd1 vssd1 vccd1 vccd1 _1779_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1701_ _2475_/Q _1706_/A _1704_/B _2476_/Q vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__a31o_1
X_2750_ _2750_/A _2048_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_2681_ _2681_/A _1965_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
X_1563_ _1634_/B _1563_/B vssd1 vssd1 vccd1 vccd1 _1611_/C sky130_fd_sc_hd__and2_1
X_1632_ _1632_/A vssd1 vssd1 vccd1 vccd1 _1639_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1498_/S _1497_/B vssd1 vssd1 vccd1 vccd1 _1495_/S sky130_fd_sc_hd__nand2_1
XFILLER_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2115_ _2115_/A vssd1 vssd1 vccd1 vccd1 _2320_/A sky130_fd_sc_hd__clkbuf_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ _2048_/A vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2733_ _2733_/A _2028_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1615_ _1577_/B _1611_/C _1611_/A vssd1 vssd1 vccd1 vccd1 _1616_/C sky130_fd_sc_hd__a21o_1
X_1546_ _1546_/A vssd1 vssd1 vccd1 vccd1 _2510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2579__7 vssd1 vssd1 vccd1 vccd1 _2579__7/HI _2683_/A sky130_fd_sc_hd__conb_1
X_1477_ _2519_/Q vssd1 vssd1 vccd1 vccd1 _1483_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2029_ _2029_/A vssd1 vssd1 vccd1 vccd1 _2029_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1331_ _2441_/Q _2440_/Q _2439_/Q _2438_/Q vssd1 vssd1 vccd1 vccd1 _1333_/C sky130_fd_sc_hd__or4_1
X_2380_ _2380_/A vssd1 vssd1 vccd1 vccd1 _2566_/D sky130_fd_sc_hd__clkbuf_1
X_1400_ _1492_/B _1584_/A vssd1 vssd1 vccd1 vccd1 _1444_/A sky130_fd_sc_hd__nor2_1
X_1262_ _2540_/Q _2539_/Q _2514_/Q _2513_/Q vssd1 vssd1 vccd1 vccd1 _1672_/A sky130_fd_sc_hd__or4_1
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2716_ _2716_/A _2008_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1529_ _2500_/Q vssd1 vssd1 vccd1 vccd1 _1591_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1880_ _1880_/A vssd1 vssd1 vccd1 vccd1 _2435_/D sky130_fd_sc_hd__clkbuf_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2501_ _2522_/CLK _2501_/D _2239_/Y vssd1 vssd1 vccd1 vccd1 _2501_/Q sky130_fd_sc_hd__dfrtp_1
X_2432_ _2439_/CLK _2432_/D _2153_/Y vssd1 vssd1 vccd1 vccd1 _2432_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2363_ _1878_/A _2382_/D _2352_/A _2381_/A vssd1 vssd1 vccd1 vccd1 _2365_/A sky130_fd_sc_hd__o211a_1
X_2294_ _2294_/A vssd1 vssd1 vccd1 vccd1 _2545_/D sky130_fd_sc_hd__clkbuf_1
X_1314_ _2570_/Q _2569_/Q _2572_/Q _2571_/Q vssd1 vssd1 vccd1 vccd1 _1318_/B sky130_fd_sc_hd__or4_1
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2655__83 vssd1 vssd1 vccd1 vccd1 _2655__83/HI _2763_/A sky130_fd_sc_hd__conb_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1932_ _1932_/A vssd1 vssd1 vccd1 vccd1 _2421_/D sky130_fd_sc_hd__clkbuf_1
X_1863_ _1866_/A _1868_/A _1928_/A vssd1 vssd1 vccd1 vccd1 _1863_/Y sky130_fd_sc_hd__a21oi_1
X_1794_ _1798_/A _1800_/A vssd1 vssd1 vccd1 vccd1 _1794_/Y sky130_fd_sc_hd__nand2_1
X_2415_ _2491_/CLK _2415_/D _2132_/Y vssd1 vssd1 vccd1 vccd1 _2415_/Q sky130_fd_sc_hd__dfrtp_1
X_2346_ _2298_/X _2343_/X _2345_/Y _2320_/X _2557_/Q vssd1 vssd1 vccd1 vccd1 _2557_/D
+ sky130_fd_sc_hd__a32o_1
X_2277_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2282_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2200_ _2202_/A vssd1 vssd1 vccd1 vccd1 _2200_/Y sky130_fd_sc_hd__inv_2
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _2134_/A vssd1 vssd1 vccd1 vccd1 _2131_/Y sky130_fd_sc_hd__inv_2
X_2062_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__inv_2
X_2625__53 vssd1 vssd1 vccd1 vccd1 _2625__53/HI _2733_/A sky130_fd_sc_hd__conb_1
X_1915_ _1915_/A vssd1 vssd1 vccd1 vccd1 _2426_/D sky130_fd_sc_hd__clkbuf_1
X_1846_ _1844_/X _2442_/Q _1840_/Y _1845_/X vssd1 vssd1 vccd1 vccd1 _2442_/D sky130_fd_sc_hd__a22o_1
X_1777_ _1777_/A _1777_/B vssd1 vssd1 vccd1 vccd1 _1781_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2329_ _2358_/B vssd1 vssd1 vccd1 vccd1 _2356_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2680_ _2680_/A _1964_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
X_1700_ _2475_/Q _1704_/B _1706_/A vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__a21boi_1
X_1631_ _2483_/Q _1646_/B vssd1 vssd1 vccd1 vccd1 _1632_/A sky130_fd_sc_hd__and2_1
X_1562_ _2487_/Q _1646_/B _1562_/C vssd1 vssd1 vccd1 vccd1 _1634_/B sky130_fd_sc_hd__and3_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1493_/A _1493_/B vssd1 vssd1 vccd1 vccd1 _1497_/B sky130_fd_sc_hd__and2_1
X_2045_ _2048_/A vssd1 vssd1 vccd1 vccd1 _2045_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2114_ _2114_/A input2/X _2323_/C vssd1 vssd1 vccd1 vccd1 _2115_/A sky130_fd_sc_hd__or3b_2
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1829_ _2417_/Q _2416_/Q vssd1 vssd1 vccd1 vccd1 _1936_/C sky130_fd_sc_hd__and2_1
XFILLER_38_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2732_ _2732_/A _2027_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
X_1614_ _1610_/Y _1616_/B _1613_/X vssd1 vssd1 vccd1 vccd1 _2493_/D sky130_fd_sc_hd__a21oi_1
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1545_ _1643_/A _1545_/B _1545_/C vssd1 vssd1 vccd1 vccd1 _1546_/A sky130_fd_sc_hd__and3_1
XFILLER_5_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1476_ _1476_/A _1476_/B vssd1 vssd1 vccd1 vccd1 _2522_/D sky130_fd_sc_hd__nor2_1
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2028_ _2029_/A vssd1 vssd1 vccd1 vccd1 _2028_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1330_ _2428_/Q _2423_/Q _2422_/Q _2429_/Q vssd1 vssd1 vccd1 vccd1 _1339_/B sky130_fd_sc_hd__or4b_2
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1261_ _1468_/A vssd1 vssd1 vccd1 vccd1 _1501_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2581__9 vssd1 vssd1 vccd1 vccd1 _2581__9/HI _2685_/A sky130_fd_sc_hd__conb_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2715_ _2715_/A _2007_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
X_1459_ _1459_/A _1459_/B vssd1 vssd1 vccd1 vccd1 _1459_/X sky130_fd_sc_hd__or2_1
X_1528_ _2499_/Q _2498_/Q _1593_/B vssd1 vssd1 vccd1 vccd1 _1559_/A sky130_fd_sc_hd__and3_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2586__14 vssd1 vssd1 vccd1 vccd1 _2586__14/HI _2690_/A sky130_fd_sc_hd__conb_1
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2431_ _2431_/CLK _2431_/D _2152_/Y vssd1 vssd1 vccd1 vccd1 _2431_/Q sky130_fd_sc_hd__dfrtp_1
X_2500_ _2522_/CLK _2500_/D _2238_/Y vssd1 vssd1 vccd1 vccd1 _2500_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2362_ _2562_/Q vssd1 vssd1 vccd1 vccd1 _2381_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2293_ _2372_/B _2320_/A _2301_/B vssd1 vssd1 vccd1 vccd1 _2294_/A sky130_fd_sc_hd__mux2_1
X_1313_ _2566_/Q _2565_/Q _2568_/Q _2567_/Q vssd1 vssd1 vccd1 vccd1 _1318_/A sky130_fd_sc_hd__or4_1
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2670__98 vssd1 vssd1 vccd1 vccd1 _2670__98/HI _2778_/A sky130_fd_sc_hd__conb_1
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1793_ _2454_/Q vssd1 vssd1 vccd1 vccd1 _1793_/Y sky130_fd_sc_hd__inv_2
X_1931_ _1928_/Y _1930_/X _2421_/Q vssd1 vssd1 vccd1 vccd1 _1932_/A sky130_fd_sc_hd__mux2_1
X_1862_ _2437_/Q _2436_/Q _1871_/B vssd1 vssd1 vccd1 vccd1 _1868_/A sky130_fd_sc_hd__and3_1
X_2414_ _2491_/CLK _2414_/D _2131_/Y vssd1 vssd1 vccd1 vccd1 _2414_/Q sky130_fd_sc_hd__dfrtp_1
X_2345_ _2350_/C vssd1 vssd1 vccd1 vccd1 _2345_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2276_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2276_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2061_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2066_/A sky130_fd_sc_hd__buf_8
X_2130_ _2134_/A vssd1 vssd1 vccd1 vccd1 _2130_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1914_ _1914_/A _1914_/B vssd1 vssd1 vccd1 vccd1 _1915_/A sky130_fd_sc_hd__and2_1
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640__68 vssd1 vssd1 vccd1 vccd1 _2640__68/HI _2748_/A sky130_fd_sc_hd__conb_1
X_1776_ _2459_/Q _1773_/A _1775_/X _1848_/A vssd1 vssd1 vccd1 vccd1 _1777_/B sky130_fd_sc_hd__a31o_1
X_1845_ _2442_/Q _1845_/B vssd1 vssd1 vccd1 vccd1 _1845_/X sky130_fd_sc_hd__or2_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2328_ _2553_/Q vssd1 vssd1 vccd1 vccd1 _2336_/B sky130_fd_sc_hd__clkbuf_1
X_2259_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2264_/A sky130_fd_sc_hd__buf_2
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ _2486_/Q _1638_/A _1639_/A vssd1 vssd1 vccd1 vccd1 _1633_/B sky130_fd_sc_hd__and3_1
X_1561_ _2494_/Q _2493_/Q _1611_/A vssd1 vssd1 vccd1 vccd1 _1564_/B sky130_fd_sc_hd__and3_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _2514_/Q _1492_/B _1501_/B vssd1 vssd1 vccd1 vccd1 _1493_/B sky130_fd_sc_hd__and3_1
X_2044_ _2048_/A vssd1 vssd1 vccd1 vccd1 _2044_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2113_ _2113_/A _2113_/B _2113_/C vssd1 vssd1 vccd1 vccd1 _2323_/C sky130_fd_sc_hd__nand3_1
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1759_ _2463_/Q _1765_/A _1765_/B _2464_/Q vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__a31o_1
X_1828_ _2415_/Q _1953_/A _2413_/Q _2412_/Q vssd1 vssd1 vccd1 vccd1 _1857_/A sky130_fd_sc_hd__and4_1
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2731_ _2731_/A _2026_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610__38 vssd1 vssd1 vccd1 vccd1 _2610__38/HI _2714_/A sky130_fd_sc_hd__conb_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_1544_ _2510_/Q _1654_/C _1544_/C vssd1 vssd1 vccd1 vccd1 _1545_/C sky130_fd_sc_hd__nand3_1
X_1613_ _1474_/X _1606_/X _1634_/A vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1475_ _2522_/Q _1650_/A _1473_/Y _1474_/X vssd1 vssd1 vccd1 vccd1 _1476_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2027_ _2029_/A vssd1 vssd1 vccd1 vccd1 _2027_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1260_ _1492_/B vssd1 vssd1 vccd1 vccd1 _1468_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2714_ _2714_/A _2004_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1527_ _2497_/Q _2496_/Q vssd1 vssd1 vccd1 vccd1 _1593_/B sky130_fd_sc_hd__and2_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1389_ _1474_/A vssd1 vssd1 vccd1 vccd1 _1555_/B sky130_fd_sc_hd__buf_2
X_1458_ _1457_/A _1457_/C _1416_/A vssd1 vssd1 vccd1 vccd1 _1459_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2430_ _2431_/CLK _2430_/D _2151_/Y vssd1 vssd1 vccd1 vccd1 _2430_/Q sky130_fd_sc_hd__dfrtp_1
X_2361_ _2302_/X _2357_/X _2360_/Y _2320_/X _2561_/Q vssd1 vssd1 vccd1 vccd1 _2561_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1312_ _1278_/X _1289_/X _2114_/A _2323_/B vssd1 vssd1 vccd1 vccd1 _1312_/Y sky130_fd_sc_hd__o211ai_1
X_2292_ _2545_/Q vssd1 vssd1 vccd1 vccd1 _2301_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2559_ _2559_/CLK _2559_/D vssd1 vssd1 vccd1 vccd1 _2559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2646__74 vssd1 vssd1 vccd1 vccd1 _2646__74/HI _2754_/A sky130_fd_sc_hd__conb_1
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1930_ _1847_/B _1928_/B _2333_/A vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__a21o_1
X_1792_ _1788_/B _1791_/Y _1787_/A _1676_/X vssd1 vssd1 vccd1 vccd1 _2455_/D sky130_fd_sc_hd__a2bb2o_1
X_1861_ _1861_/A _1933_/A _1875_/B _1861_/D vssd1 vssd1 vccd1 vccd1 _1871_/B sky130_fd_sc_hd__and4_1
X_2413_ _2491_/CLK _2413_/D _2130_/Y vssd1 vssd1 vccd1 vccd1 _2413_/Q sky130_fd_sc_hd__dfrtp_1
X_2344_ _2556_/Q _2557_/Q _2344_/C vssd1 vssd1 vccd1 vccd1 _2350_/C sky130_fd_sc_hd__and3_1
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2275_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2275_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2060_ _2060_/A vssd1 vssd1 vccd1 vccd1 _2060_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _2425_/Q _1885_/A _1916_/B _2426_/Q vssd1 vssd1 vccd1 vccd1 _1914_/B sky130_fd_sc_hd__a31o_1
X_1775_ _1785_/A _1788_/A _1787_/A _1787_/B vssd1 vssd1 vccd1 vccd1 _1775_/X sky130_fd_sc_hd__and4_1
X_1844_ _1903_/A vssd1 vssd1 vccd1 vccd1 _1844_/X sky130_fd_sc_hd__clkbuf_2
X_2327_ _2327_/A _2327_/B vssd1 vssd1 vccd1 vccd1 _2552_/D sky130_fd_sc_hd__nor2_1
X_2258_ _2258_/A vssd1 vssd1 vccd1 vccd1 _2258_/Y sky130_fd_sc_hd__inv_2
X_2189_ _2190_/A vssd1 vssd1 vccd1 vccd1 _2189_/Y sky130_fd_sc_hd__inv_2
X_2616__44 vssd1 vssd1 vccd1 vccd1 _2616__44/HI _2720_/A sky130_fd_sc_hd__conb_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2560_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1560_ _2502_/Q _2501_/Q _1591_/S _1589_/B vssd1 vssd1 vccd1 vccd1 _1580_/A sky130_fd_sc_hd__and4_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2112_ _2572_/Q _2410_/Q _2112_/C _2119_/A vssd1 vssd1 vccd1 vccd1 _2126_/B sky130_fd_sc_hd__nand4_1
X_1491_ _2513_/Q _1509_/A _1511_/S vssd1 vssd1 vccd1 vccd1 _1501_/B sky130_fd_sc_hd__and3_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2043_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2048_/A sky130_fd_sc_hd__buf_6
X_1827_ _2414_/Q vssd1 vssd1 vccd1 vccd1 _1953_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1758_ _2461_/Q _1800_/A _1758_/C vssd1 vssd1 vccd1 vccd1 _1765_/B sky130_fd_sc_hd__and3_1
X_1689_ _2459_/Q _2454_/Q _1798_/A vssd1 vssd1 vccd1 vccd1 _1690_/C sky130_fd_sc_hd__and3_1
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ _2730_/A _2025_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
X_1543_ _1612_/A vssd1 vssd1 vccd1 vccd1 _1654_/C sky130_fd_sc_hd__clkbuf_2
X_1612_ _1612_/A vssd1 vssd1 vccd1 vccd1 _1634_/A sky130_fd_sc_hd__clkbuf_2
X_1474_ _1474_/A vssd1 vssd1 vccd1 vccd1 _1474_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2026_ _2029_/A vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2713_ _2713_/A _2003_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1526_ _2506_/Q _2505_/Q _1578_/S _2503_/Q vssd1 vssd1 vccd1 vccd1 _1567_/A sky130_fd_sc_hd__and4_1
X_1457_ _1457_/A _1457_/B _1457_/C vssd1 vssd1 vccd1 vccd1 _1457_/X sky130_fd_sc_hd__and3_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1388_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1474_/A sky130_fd_sc_hd__clkbuf_2
X_2009_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2009_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1311_ input2/X vssd1 vssd1 vccd1 vccd1 _2323_/B sky130_fd_sc_hd__inv_2
X_2360_ _2382_/D vssd1 vssd1 vccd1 vccd1 _2360_/Y sky130_fd_sc_hd__inv_2
X_2291_ _2399_/A vssd1 vssd1 vccd1 vccd1 _2372_/B sky130_fd_sc_hd__buf_2
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2558_ _2559_/CLK _2558_/D vssd1 vssd1 vccd1 vccd1 _2558_/Q sky130_fd_sc_hd__dfxtp_1
X_2489_ _2506_/CLK _2489_/D _2224_/Y vssd1 vssd1 vccd1 vccd1 _2489_/Q sky130_fd_sc_hd__dfrtp_1
X_1509_ _1509_/A _1511_/S vssd1 vssd1 vccd1 vccd1 _1509_/X sky130_fd_sc_hd__or2_1
X_2661__89 vssd1 vssd1 vccd1 vccd1 _2661__89/HI _2769_/A sky130_fd_sc_hd__conb_1
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ _1925_/A _1874_/B _1923_/B vssd1 vssd1 vccd1 vccd1 _1861_/D sky130_fd_sc_hd__and3_1
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1791_ _1787_/A _1787_/B _1706_/A vssd1 vssd1 vccd1 vccd1 _1791_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2412_ _2544_/CLK _2412_/D _2323_/B vssd1 vssd1 vccd1 vccd1 _2412_/Q sky130_fd_sc_hd__dfrtp_1
X_2343_ _2356_/A _2109_/C _2557_/Q vssd1 vssd1 vccd1 vccd1 _2343_/X sky130_fd_sc_hd__a21o_1
X_2274_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2274_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1989_ _1992_/A vssd1 vssd1 vccd1 vccd1 _1989_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ _2427_/Q _1914_/A _1911_/Y _1909_/X vssd1 vssd1 vccd1 vccd1 _2427_/D sky130_fd_sc_hd__a22o_1
X_1843_ _2333_/A vssd1 vssd1 vccd1 vccd1 _1903_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1774_ _2459_/Q _1774_/B _1774_/C vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__and3_1
X_2326_ _1795_/X _2318_/A _2352_/A _2552_/Q vssd1 vssd1 vccd1 vccd1 _2327_/B sky130_fd_sc_hd__o211a_1
X_2257_ _2258_/A vssd1 vssd1 vccd1 vccd1 _2257_/Y sky130_fd_sc_hd__inv_2
X_2188_ _2190_/A vssd1 vssd1 vccd1 vccd1 _2188_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2631__59 vssd1 vssd1 vccd1 vccd1 _2631__59/HI _2739_/A sky130_fd_sc_hd__conb_1
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1670_/D _1513_/A vssd1 vssd1 vccd1 vccd1 _1490_/Y sky130_fd_sc_hd__nand2_1
X_2111_ _2111_/A _2393_/B vssd1 vssd1 vccd1 vccd1 _2119_/A sky130_fd_sc_hd__nor2_1
X_2042_ _2042_/A vssd1 vssd1 vccd1 vccd1 _2042_/Y sky130_fd_sc_hd__inv_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1826_ _2438_/Q vssd1 vssd1 vccd1 vccd1 _1866_/A sky130_fd_sc_hd__clkbuf_1
X_1757_ _1757_/A vssd1 vssd1 vccd1 vccd1 _1757_/Y sky130_fd_sc_hd__inv_2
X_1688_ _2453_/Q vssd1 vssd1 vccd1 vccd1 _1798_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2309_ _2549_/Q vssd1 vssd1 vccd1 vccd1 _2314_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1611_ _1611_/A _1639_/B _1611_/C vssd1 vssd1 vccd1 vccd1 _1616_/B sky130_fd_sc_hd__nand3_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1542_ _1639_/B _1544_/C _2510_/Q vssd1 vssd1 vccd1 vccd1 _1545_/B sky130_fd_sc_hd__a21o_1
X_1473_ _1473_/A vssd1 vssd1 vccd1 vccd1 _1473_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2025_ _2029_/A vssd1 vssd1 vccd1 vccd1 _2025_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1809_ _1806_/B _1808_/X _2450_/Q _1703_/X vssd1 vssd1 vccd1 vccd1 _2450_/D sky130_fd_sc_hd__a2bb2o_1
X_2601__29 vssd1 vssd1 vccd1 vccd1 _2601__29/HI _2705_/A sky130_fd_sc_hd__conb_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2667__95 vssd1 vssd1 vccd1 vccd1 _2667__95/HI _2775_/A sky130_fd_sc_hd__conb_1
XFILLER_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2712_/A _2002_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
X_2574_ _2574_/CLK _2574_/D vssd1 vssd1 vccd1 vccd1 _2574_/Q sky130_fd_sc_hd__dfxtp_1
X_1387_ _1387_/A _1387_/B vssd1 vssd1 vccd1 vccd1 _1415_/A sky130_fd_sc_hd__nand2_1
X_1525_ _2504_/Q vssd1 vssd1 vccd1 vccd1 _1578_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_1456_ _1465_/A _1467_/A _1472_/D _1468_/C vssd1 vssd1 vccd1 vccd1 _1457_/C sky130_fd_sc_hd__and4_1
X_2008_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1310_ _1387_/A vssd1 vssd1 vccd1 vccd1 _2114_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2290_ _2290_/A vssd1 vssd1 vccd1 vccd1 _2290_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2557_ _2560_/CLK _2557_/D vssd1 vssd1 vccd1 vccd1 _2557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ _2506_/CLK _2488_/D _2223_/Y vssd1 vssd1 vccd1 vccd1 _2488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1439_ _1445_/S _1442_/A _1442_/B vssd1 vssd1 vccd1 vccd1 _1439_/X sky130_fd_sc_hd__and3_1
X_1508_ _1508_/A vssd1 vssd1 vccd1 vccd1 _2513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2637__65 vssd1 vssd1 vccd1 vccd1 _2637__65/HI _2745_/A sky130_fd_sc_hd__conb_1
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1790_ _1788_/A _1761_/X _1708_/A _1789_/Y vssd1 vssd1 vccd1 vccd1 _2456_/D sky130_fd_sc_hd__a22o_1
X_2411_ _2574_/CLK _2411_/D vssd1 vssd1 vccd1 vccd1 _2411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2342_ _2342_/A _2342_/B vssd1 vssd1 vccd1 vccd1 _2556_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2273_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2273_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1988_ _1992_/A vssd1 vssd1 vccd1 vccd1 _1988_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1911_ _2427_/Q _1911_/B vssd1 vssd1 vccd1 vccd1 _1911_/Y sky130_fd_sc_hd__nor2_1
X_1773_ _1773_/A _1785_/A _1789_/A vssd1 vssd1 vccd1 vccd1 _1774_/C sky130_fd_sc_hd__and3_1
X_1842_ _1824_/X _1825_/Y _1840_/Y _1841_/X vssd1 vssd1 vccd1 vccd1 _2443_/D sky130_fd_sc_hd__o31a_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2187_ _2190_/A vssd1 vssd1 vccd1 vccd1 _2187_/Y sky130_fd_sc_hd__inv_2
X_2325_ _2403_/A vssd1 vssd1 vccd1 vccd1 _2352_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2256_ _2258_/A vssd1 vssd1 vccd1 vccd1 _2256_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2607__35 vssd1 vssd1 vccd1 vccd1 _2607__35/HI _2711_/A sky130_fd_sc_hd__conb_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2041_ _2042_/A vssd1 vssd1 vccd1 vccd1 _2041_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2110_ _2569_/Q _2110_/B _2358_/B _2358_/C vssd1 vssd1 vccd1 vccd1 _2393_/B sky130_fd_sc_hd__nand4_1
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1756_ _1734_/X _1753_/Y _1754_/X _1755_/X _1754_/A vssd1 vssd1 vccd1 vccd1 _2465_/D
+ sky130_fd_sc_hd__a32o_1
X_1825_ _2443_/Q vssd1 vssd1 vccd1 vccd1 _1825_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1687_ _2458_/Q _1785_/A _1788_/A _2455_/Q vssd1 vssd1 vccd1 vccd1 _1690_/B sky130_fd_sc_hd__and4_1
X_2308_ _2306_/Y _2302_/X _2307_/X _2299_/X _2548_/Q vssd1 vssd1 vccd1 vccd1 _2548_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2239_ _2240_/A vssd1 vssd1 vccd1 vccd1 _2239_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1610_ _2493_/Q vssd1 vssd1 vccd1 vccd1 _1610_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1541_ _2509_/Q _2508_/Q _2507_/Q _1553_/B vssd1 vssd1 vccd1 vccd1 _1544_/C sky130_fd_sc_hd__and4_1
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1472_ _1472_/A _1480_/A _2519_/Q _1472_/D vssd1 vssd1 vccd1 vccd1 _1473_/A sky130_fd_sc_hd__and4_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2024_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2029_/A sky130_fd_sc_hd__buf_8
XFILLER_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2598__26 vssd1 vssd1 vccd1 vccd1 _2598__26/HI _2702_/A sky130_fd_sc_hd__conb_1
X_1808_ _1803_/A _1803_/B _1737_/B _1795_/X vssd1 vssd1 vccd1 vccd1 _1808_/X sky130_fd_sc_hd__a211o_1
X_1739_ _2465_/Q vssd1 vssd1 vccd1 vccd1 _1754_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2711_ _2711_/A _2093_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
X_1524_ _1612_/A vssd1 vssd1 vccd1 vccd1 _1639_/B sky130_fd_sc_hd__clkbuf_2
X_2573_ _2574_/CLK _2573_/D vssd1 vssd1 vccd1 vccd1 _2573_/Q sky130_fd_sc_hd__dfxtp_1
X_2675__103 vssd1 vssd1 vccd1 vccd1 _2675__103/HI _2783_/A sky130_fd_sc_hd__conb_1
X_1386_ _1386_/A vssd1 vssd1 vccd1 vccd1 _2539_/D sky130_fd_sc_hd__inv_2
X_1455_ _1455_/A _1455_/B vssd1 vssd1 vccd1 vccd1 _1472_/D sky130_fd_sc_hd__and2_1
X_2007_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2007_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2556_ _2560_/CLK _2556_/D vssd1 vssd1 vccd1 vccd1 _2556_/Q sky130_fd_sc_hd__dfxtp_1
X_2487_ _2491_/CLK _2487_/D _2221_/Y vssd1 vssd1 vccd1 vccd1 _2487_/Q sky130_fd_sc_hd__dfrtp_1
X_1507_ _1507_/A _1507_/B vssd1 vssd1 vccd1 vccd1 _1508_/A sky130_fd_sc_hd__and2_1
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1369_ _1387_/B vssd1 vssd1 vccd1 vccd1 _2113_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1438_ _1492_/B _1438_/B _1453_/B vssd1 vssd1 vccd1 vccd1 _1442_/B sky130_fd_sc_hd__and3_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2582__10 vssd1 vssd1 vccd1 vccd1 _2582__10/HI _2686_/A sky130_fd_sc_hd__conb_1
XFILLER_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2341_ _1795_/X _2344_/C _2352_/A _2556_/Q vssd1 vssd1 vccd1 vccd1 _2342_/B sky130_fd_sc_hd__o211a_1
X_2410_ _2574_/CLK _2410_/D vssd1 vssd1 vccd1 vccd1 _2410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2272_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2272_/Y sky130_fd_sc_hd__inv_2
X_1987_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1992_/A sky130_fd_sc_hd__buf_8
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2539_ _2572_/CLK _2539_/D _2285_/Y vssd1 vssd1 vccd1 vccd1 _2539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1910_ _1911_/B _1909_/X _1878_/A vssd1 vssd1 vccd1 vccd1 _1914_/A sky130_fd_sc_hd__o21ai_1
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1772_ _1788_/A _1787_/A _1787_/B vssd1 vssd1 vccd1 vccd1 _1789_/A sky130_fd_sc_hd__and3_1
X_1841_ _2442_/Q _1821_/X _1845_/B _2443_/Q vssd1 vssd1 vccd1 vccd1 _1841_/X sky130_fd_sc_hd__a31o_1
XFILLER_8_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2324_ _2324_/A vssd1 vssd1 vccd1 vccd1 _2403_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2186_ _2190_/A vssd1 vssd1 vccd1 vccd1 _2186_/Y sky130_fd_sc_hd__inv_2
X_2255_ _2258_/A vssd1 vssd1 vccd1 vccd1 _2255_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _2042_/A vssd1 vssd1 vccd1 vccd1 _2040_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1755_ _1761_/A vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__clkbuf_2
X_1686_ _2456_/Q vssd1 vssd1 vccd1 vccd1 _1788_/A sky130_fd_sc_hd__clkbuf_1
X_1824_ _2333_/A vssd1 vssd1 vccd1 vccd1 _1824_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2307_ _2301_/A _2301_/B _2301_/C _2548_/Q vssd1 vssd1 vccd1 vccd1 _2307_/X sky130_fd_sc_hd__a31o_1
X_2238_ _2240_/A vssd1 vssd1 vccd1 vccd1 _2238_/Y sky130_fd_sc_hd__inv_2
X_2169_ _2171_/A vssd1 vssd1 vccd1 vccd1 _2169_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1540_ _1567_/A _1570_/B vssd1 vssd1 vccd1 vccd1 _1553_/B sky130_fd_sc_hd__and2_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1471_ _2520_/Q vssd1 vssd1 vccd1 vccd1 _1480_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2023_ _2023_/A vssd1 vssd1 vccd1 vccd1 _2023_/Y sky130_fd_sc_hd__inv_2
X_1807_ _2451_/Q _1761_/X _1715_/X _1806_/X vssd1 vssd1 vccd1 vccd1 _2451_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1738_ _1734_/X _1732_/B _1736_/X _1737_/X vssd1 vssd1 vccd1 vccd1 _2469_/D sky130_fd_sc_hd__a31o_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2568_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_1669_ _1669_/A _1669_/B _1669_/C _1669_/D vssd1 vssd1 vccd1 vccd1 _1669_/X sky130_fd_sc_hd__or4_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ _2710_/A _2001_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1523_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1612_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2572_ _2572_/CLK _2572_/D vssd1 vssd1 vccd1 vccd1 _2572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1454_ _1451_/X _1452_/Y _1453_/X _1402_/X _1453_/A vssd1 vssd1 vccd1 vccd1 _2527_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1385_ _1383_/Y _2539_/Q _1385_/S vssd1 vssd1 vccd1 vccd1 _1386_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2006_ _2030_/A vssd1 vssd1 vccd1 vccd1 _2011_/A sky130_fd_sc_hd__buf_8
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2658__86 vssd1 vssd1 vccd1 vccd1 _2658__86/HI _2766_/A sky130_fd_sc_hd__conb_1
XFILLER_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2555_ _2560_/CLK _2555_/D vssd1 vssd1 vccd1 vccd1 _2555_/Q sky130_fd_sc_hd__dfxtp_1
X_2486_ _2491_/CLK _2486_/D _2220_/Y vssd1 vssd1 vccd1 vccd1 _2486_/Q sky130_fd_sc_hd__dfrtp_1
X_1506_ _1474_/A _1505_/Y _1382_/A _2513_/Q vssd1 vssd1 vccd1 vccd1 _1507_/B sky130_fd_sc_hd__a2bb2o_1
X_1437_ _2532_/Q _2531_/Q vssd1 vssd1 vccd1 vccd1 _1437_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1299_ _2492_/Q _2491_/Q _2490_/Q _2489_/Q vssd1 vssd1 vccd1 vccd1 _1303_/A sky130_fd_sc_hd__or4_1
X_1368_ _2541_/Q _2540_/Q _1375_/B vssd1 vssd1 vccd1 vccd1 _1372_/B sky130_fd_sc_hd__and3_1
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _2372_/B _2344_/C _2556_/Q vssd1 vssd1 vccd1 vccd1 _2342_/A sky130_fd_sc_hd__a21oi_1
X_2271_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2276_/A sky130_fd_sc_hd__buf_2
X_2628__56 vssd1 vssd1 vccd1 vccd1 _2628__56/HI _2736_/A sky130_fd_sc_hd__conb_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1986_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1986_/Y sky130_fd_sc_hd__inv_2
X_2469_ _2559_/CLK _2469_/D _2199_/Y vssd1 vssd1 vccd1 vccd1 _2469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2538_ _2568_/CLK _2538_/D _2284_/Y vssd1 vssd1 vccd1 vccd1 _2538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2642__70 vssd1 vssd1 vccd1 vccd1 _2642__70/HI _2750_/A sky130_fd_sc_hd__conb_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1840_ _2442_/Q _1845_/B _1947_/A vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1771_ _2454_/Q _1798_/A _1771_/C vssd1 vssd1 vccd1 vccd1 _1787_/B sky130_fd_sc_hd__and3_1
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2323_ _1387_/A _2323_/B _2323_/C vssd1 vssd1 vccd1 vccd1 _2324_/A sky130_fd_sc_hd__and3b_1
X_2254_ _2258_/A vssd1 vssd1 vccd1 vccd1 _2254_/Y sky130_fd_sc_hd__inv_2
X_2185_ _2197_/A vssd1 vssd1 vccd1 vccd1 _2190_/A sky130_fd_sc_hd__buf_2
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ _1973_/A vssd1 vssd1 vccd1 vccd1 _1969_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1823_ _2725_/A _1822_/X _1712_/C vssd1 vssd1 vccd1 vccd1 _2444_/D sky130_fd_sc_hd__a21o_1
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1754_ _1754_/A _1757_/A vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__or2_1
X_1685_ _2457_/Q vssd1 vssd1 vccd1 vccd1 _1785_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2306_ _2314_/B vssd1 vssd1 vccd1 vccd1 _2306_/Y sky130_fd_sc_hd__inv_2
X_2237_ _2240_/A vssd1 vssd1 vccd1 vccd1 _2237_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _2171_/A vssd1 vssd1 vccd1 vccd1 _2168_/Y sky130_fd_sc_hd__inv_2
X_2099_ _2564_/Q vssd1 vssd1 vccd1 vccd1 _2382_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2612__40 vssd1 vssd1 vccd1 vccd1 _2612__40/HI _2716_/A sky130_fd_sc_hd__conb_1
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1470_ _1470_/A vssd1 vssd1 vccd1 vccd1 _2523_/D sky130_fd_sc_hd__inv_2
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2022_ _2023_/A vssd1 vssd1 vccd1 vccd1 _2022_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1806_ _2451_/Q _1806_/B vssd1 vssd1 vccd1 vccd1 _1806_/X sky130_fd_sc_hd__xor2_1
X_2786_ _2786_/A _2091_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1737_ _2469_/Q _1737_/B vssd1 vssd1 vccd1 vccd1 _1737_/X sky130_fd_sc_hd__and2_1
X_1599_ _1474_/X _1593_/B _1593_/C _1657_/A vssd1 vssd1 vccd1 vccd1 _1600_/B sky130_fd_sc_hd__o22a_1
X_1668_ _1668_/A _1668_/B _1435_/A _2533_/Q vssd1 vssd1 vccd1 vccd1 _1669_/D sky130_fd_sc_hd__or4bb_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2589__17 vssd1 vssd1 vccd1 vccd1 _2589__17/HI _2693_/A sky130_fd_sc_hd__conb_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1522_ _1416_/A _1658_/B _1521_/Y vssd1 vssd1 vccd1 vccd1 _1549_/A sky130_fd_sc_hd__o21a_1
X_2571_ _2572_/CLK _2571_/D vssd1 vssd1 vccd1 vccd1 _2571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1453_ _1453_/A _1453_/B vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__or2_1
X_2005_ input1/X vssd1 vssd1 vccd1 vccd1 _2030_/A sky130_fd_sc_hd__buf_2
X_1384_ _1468_/A _1384_/B _1420_/B vssd1 vssd1 vccd1 vccd1 _1385_/S sky130_fd_sc_hd__and3_1
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2769_ _2769_/A _2071_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2554_ _2574_/CLK _2554_/D vssd1 vssd1 vccd1 vccd1 _2554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2485_ _2491_/CLK _2485_/D _2219_/Y vssd1 vssd1 vccd1 vccd1 _2485_/Q sky130_fd_sc_hd__dfrtp_1
X_1505_ _1509_/A _1511_/S vssd1 vssd1 vccd1 vccd1 _1505_/Y sky130_fd_sc_hd__nand2_1
X_1436_ _1457_/B _1435_/Y _1459_/A vssd1 vssd1 vccd1 vccd1 _1436_/X sky130_fd_sc_hd__a21o_1
X_1367_ _2539_/Q _1492_/B _1384_/B _1420_/B vssd1 vssd1 vccd1 vccd1 _1375_/B sky130_fd_sc_hd__and4_1
X_1298_ _1298_/A _1298_/B _1298_/C _1298_/D vssd1 vssd1 vccd1 vccd1 _1665_/C sky130_fd_sc_hd__nor4_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2270_ _2270_/A vssd1 vssd1 vccd1 vccd1 _2270_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1985_/Y sky130_fd_sc_hd__inv_2
X_2537_ _2537_/CLK _2537_/D _2282_/Y vssd1 vssd1 vccd1 vccd1 _2537_/Q sky130_fd_sc_hd__dfrtp_1
X_2468_ _2559_/CLK _2468_/D _2198_/Y vssd1 vssd1 vccd1 vccd1 _2468_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2399_ _2399_/A _2407_/D vssd1 vssd1 vccd1 vccd1 _2399_/X sky130_fd_sc_hd__and2_1
X_1419_ _1419_/A _1513_/A vssd1 vssd1 vccd1 vccd1 _1419_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1770_ _2455_/Q vssd1 vssd1 vccd1 vccd1 _1787_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2184_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2184_/Y sky130_fd_sc_hd__inv_2
X_2322_ _2372_/B _2318_/A _2552_/Q vssd1 vssd1 vccd1 vccd1 _2327_/A sky130_fd_sc_hd__a21oi_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2253_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2258_/A sky130_fd_sc_hd__buf_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_1899_ _1902_/A _1906_/A _1906_/B _2430_/Q vssd1 vssd1 vccd1 vccd1 _1899_/X sky130_fd_sc_hd__a31o_1
X_1968_ _2093_/A vssd1 vssd1 vccd1 vccd1 _1973_/A sky130_fd_sc_hd__buf_6
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1753_ _1754_/A _1757_/A vssd1 vssd1 vccd1 vccd1 _1753_/Y sky130_fd_sc_hd__nand2_1
X_1822_ _1821_/X _1710_/B _1658_/Y vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__a21o_1
X_1684_ _1771_/C vssd1 vssd1 vccd1 vccd1 _1800_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2167_ _2171_/A vssd1 vssd1 vccd1 vccd1 _2167_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2305_ _2305_/A vssd1 vssd1 vccd1 vccd1 _2314_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2236_ _2240_/A vssd1 vssd1 vccd1 vccd1 _2236_/Y sky130_fd_sc_hd__inv_2
X_2098_ _2566_/Q _2565_/Q _2567_/Q vssd1 vssd1 vccd1 vccd1 _2382_/B sky130_fd_sc_hd__and3_1
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2021_ _2023_/A vssd1 vssd1 vccd1 vccd1 _2021_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1805_ _1715_/A _1800_/Y _1804_/X _1680_/X _2452_/Q vssd1 vssd1 vccd1 vccd1 _2452_/D
+ sky130_fd_sc_hd__a32o_1
X_1736_ _1757_/A _1720_/C _2469_/Q vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__a21o_1
X_2785_ _2785_/A _2090_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ _1667_/A vssd1 vssd1 vccd1 vccd1 _2478_/D sky130_fd_sc_hd__clkbuf_1
X_1598_ _2496_/Q _1595_/X _2497_/Q vssd1 vssd1 vccd1 vccd1 _1600_/A sky130_fd_sc_hd__a21oi_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2219_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2219_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2570_ _2572_/CLK _2570_/D vssd1 vssd1 vccd1 vccd1 _2570_/Q sky130_fd_sc_hd__dfxtp_1
X_1521_ _1415_/A _1278_/X _1382_/A vssd1 vssd1 vccd1 vccd1 _1521_/Y sky130_fd_sc_hd__o21ai_1
X_1383_ _2539_/Q _1650_/A vssd1 vssd1 vccd1 vccd1 _1383_/Y sky130_fd_sc_hd__nand2_1
X_1452_ _1453_/A _1453_/B vssd1 vssd1 vccd1 vccd1 _1452_/Y sky130_fd_sc_hd__nand2_1
X_2004_ _2004_/A vssd1 vssd1 vccd1 vccd1 _2004_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2768_ _2768_/A _2070_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_1719_ _1771_/C _1758_/C _1719_/C vssd1 vssd1 vccd1 vccd1 _1740_/C sky130_fd_sc_hd__and3_1
X_2699_ _2699_/A _1988_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2649__77 vssd1 vssd1 vccd1 vccd1 _2649__77/HI _2757_/A sky130_fd_sc_hd__conb_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663__91 vssd1 vssd1 vccd1 vccd1 _2663__91/HI _2771_/A sky130_fd_sc_hd__conb_1
XFILLER_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2553_ _2574_/CLK _2553_/D vssd1 vssd1 vccd1 vccd1 _2553_/Q sky130_fd_sc_hd__dfxtp_1
X_1504_ _1507_/A _1503_/Y _1493_/B vssd1 vssd1 vccd1 vccd1 _2514_/D sky130_fd_sc_hd__a21oi_1
X_2484_ _2491_/CLK _2484_/D _2218_/Y vssd1 vssd1 vccd1 vccd1 _2484_/Q sky130_fd_sc_hd__dfrtp_1
X_1435_ _1435_/A _1435_/B _1453_/B vssd1 vssd1 vccd1 vccd1 _1435_/Y sky130_fd_sc_hd__nand3_1
X_1366_ _1438_/B _1425_/B _1434_/A _1393_/C vssd1 vssd1 vccd1 vccd1 _1420_/B sky130_fd_sc_hd__and4_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1297_ _2504_/Q _2503_/Q _2502_/Q _2501_/Q vssd1 vssd1 vccd1 vccd1 _1298_/D sky130_fd_sc_hd__or4_1
XFILLER_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1984_/Y sky130_fd_sc_hd__inv_2
X_2467_ _2560_/CLK _2467_/D _2196_/Y vssd1 vssd1 vccd1 vccd1 _2467_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_2536_ _2537_/CLK _2536_/D _2281_/Y vssd1 vssd1 vccd1 vccd1 _2536_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _2571_/Q _2396_/Y _2397_/X _2393_/Y vssd1 vssd1 vccd1 vccd1 _2571_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1349_ _2531_/Q vssd1 vssd1 vccd1 vccd1 _1435_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2619__47 vssd1 vssd1 vccd1 vccd1 _2619__47/HI _2723_/A sky130_fd_sc_hd__conb_1
X_1418_ _1413_/A _1402_/X _1417_/X vssd1 vssd1 vccd1 vccd1 _2536_/D sky130_fd_sc_hd__a21bo_1
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2633__61 vssd1 vssd1 vccd1 vccd1 _2633__61/HI _2741_/A sky130_fd_sc_hd__conb_1
X_2321_ _2298_/X _2318_/Y _2319_/X _2320_/X _2551_/Q vssd1 vssd1 vccd1 vccd1 _2551_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2183_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__inv_2
X_2252_ _2252_/A vssd1 vssd1 vccd1 vccd1 _2252_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1898_ _2431_/Q _1896_/X _1897_/X vssd1 vssd1 vccd1 vccd1 _2431_/D sky130_fd_sc_hd__a21bo_1
X_1967_ _1967_/A vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__inv_2
X_2519_ _2522_/CLK _2519_/D _2261_/Y vssd1 vssd1 vccd1 vccd1 _2519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1683_ _2449_/Q _1812_/A _1683_/C vssd1 vssd1 vccd1 vccd1 _1771_/C sky130_fd_sc_hd__and3_1
X_1752_ _2466_/Q _1703_/X _1715_/X _1751_/Y vssd1 vssd1 vccd1 vccd1 _2466_/D sky130_fd_sc_hd__a22o_1
X_1821_ _1847_/B vssd1 vssd1 vccd1 vccd1 _1821_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2304_ _2301_/Y _2302_/X _2303_/X _2299_/X _2301_/C vssd1 vssd1 vccd1 vccd1 _2547_/D
+ sky130_fd_sc_hd__a32o_1
X_2166_ _2166_/A vssd1 vssd1 vccd1 vccd1 _2171_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2097_ _2570_/Q _2571_/Q vssd1 vssd1 vccd1 vccd1 _2111_/A sky130_fd_sc_hd__nand2_1
X_2235_ _2259_/A vssd1 vssd1 vccd1 vccd1 _2240_/A sky130_fd_sc_hd__buf_2
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2603__31 vssd1 vssd1 vccd1 vccd1 _2603__31/HI _2707_/A sky130_fd_sc_hd__conb_1
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2020_ _2023_/A vssd1 vssd1 vccd1 vccd1 _2020_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1804_ _2451_/Q _1806_/B _2452_/Q vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__a21o_1
X_1735_ _1740_/C vssd1 vssd1 vccd1 vccd1 _1757_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1666_ _1666_/A _1666_/B vssd1 vssd1 vccd1 vccd1 _1667_/A sky130_fd_sc_hd__or2_1
X_2784_ _2784_/A _2089_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _1637_/A _1597_/B _1597_/C vssd1 vssd1 vccd1 vccd1 _2498_/D sky130_fd_sc_hd__nor3_1
X_2149_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2149_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2218_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2218_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1520_ _1413_/B _1289_/X _1519_/X _1278_/X vssd1 vssd1 vccd1 vccd1 _1658_/B sky130_fd_sc_hd__a22oi_2
X_1382_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1650_/A sky130_fd_sc_hd__clkbuf_4
X_1451_ _1457_/B vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__clkbuf_2
X_2003_ _2004_/A vssd1 vssd1 vccd1 vccd1 _2003_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2594__22 vssd1 vssd1 vccd1 vccd1 _2594__22/HI _2698_/A sky130_fd_sc_hd__conb_1
X_2767_ _2767_/A _2069_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
X_1718_ _2470_/Q vssd1 vssd1 vccd1 vccd1 _1732_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1649_ _2481_/Q _1654_/A _2479_/Q _1577_/B _2482_/Q vssd1 vssd1 vccd1 vccd1 _1650_/C
+ sky130_fd_sc_hd__a41o_1
X_2698_ _2698_/A _1986_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2537_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2552_ _2560_/CLK _2552_/D vssd1 vssd1 vccd1 vccd1 _2552_/Q sky130_fd_sc_hd__dfxtp_1
X_2483_ _2544_/CLK _2483_/D _2217_/Y vssd1 vssd1 vccd1 vccd1 _2483_/Q sky130_fd_sc_hd__dfrtp_1
X_1503_ _2514_/Q _1503_/B vssd1 vssd1 vccd1 vccd1 _1503_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1434_ _1434_/A vssd1 vssd1 vccd1 vccd1 _1453_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1365_ _1668_/A _1430_/A vssd1 vssd1 vccd1 vccd1 _1393_/C sky130_fd_sc_hd__and2_1
X_1296_ _2500_/Q _2499_/Q _2498_/Q _2497_/Q vssd1 vssd1 vccd1 vccd1 _1298_/C sky130_fd_sc_hd__or4_2
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1983_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1983_/Y sky130_fd_sc_hd__inv_2
X_2466_ _2559_/CLK _2466_/D _2195_/Y vssd1 vssd1 vccd1 vccd1 _2466_/Q sky130_fd_sc_hd__dfrtp_1
X_2577__5 vssd1 vssd1 vccd1 vccd1 _2577__5/HI _2681_/A sky130_fd_sc_hd__conb_1
X_1417_ _1417_/A _1417_/B _1658_/A vssd1 vssd1 vccd1 vccd1 _1417_/X sky130_fd_sc_hd__or3_1
X_2535_ _2572_/CLK _2535_/D _2280_/Y vssd1 vssd1 vccd1 vccd1 _2535_/Q sky130_fd_sc_hd__dfrtp_2
X_1279_ _2474_/Q _2473_/Q _2472_/Q _2471_/Q vssd1 vssd1 vccd1 vccd1 _1281_/C sky130_fd_sc_hd__or4_1
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2397_ _2571_/Q _2570_/Q vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__and2b_1
X_1348_ _2532_/Q vssd1 vssd1 vccd1 vccd1 _1668_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2320_ _2320_/A vssd1 vssd1 vccd1 vccd1 _2320_/X sky130_fd_sc_hd__clkbuf_2
X_2251_ _2252_/A vssd1 vssd1 vccd1 vccd1 _2251_/Y sky130_fd_sc_hd__inv_2
X_2182_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2182_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1966_ _1967_/A vssd1 vssd1 vccd1 vccd1 _1966_/Y sky130_fd_sc_hd__inv_2
X_1897_ _2431_/Q _1911_/B _1897_/C vssd1 vssd1 vccd1 vccd1 _1897_/X sky130_fd_sc_hd__or3_1
X_2449_ _2464_/CLK _2449_/D _2175_/Y vssd1 vssd1 vccd1 vccd1 _2449_/Q sky130_fd_sc_hd__dfrtp_1
X_2518_ _2526_/CLK _2518_/D _2260_/Y vssd1 vssd1 vccd1 vccd1 _2518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1820_ _1820_/A vssd1 vssd1 vccd1 vccd1 _2445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1682_ _2452_/Q _2451_/Q _2450_/Q vssd1 vssd1 vccd1 vccd1 _1683_/C sky130_fd_sc_hd__and3_1
X_1751_ _1751_/A _1751_/B vssd1 vssd1 vccd1 vccd1 _1751_/Y sky130_fd_sc_hd__nor2_1
X_2303_ _2301_/A _2301_/B _2301_/C vssd1 vssd1 vccd1 vccd1 _2303_/X sky130_fd_sc_hd__a21o_1
X_2234_ _2234_/A vssd1 vssd1 vccd1 vccd1 _2259_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2165_ _2165_/A vssd1 vssd1 vccd1 vccd1 _2165_/Y sky130_fd_sc_hd__inv_2
X_2096_ _2574_/Q _2573_/Q vssd1 vssd1 vccd1 vccd1 _2112_/C sky130_fd_sc_hd__and2_1
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2431_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_1949_ _2413_/Q vssd1 vssd1 vccd1 vccd1 _1956_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2783_ _2783_/A _2088_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1803_ _1803_/A _1803_/B vssd1 vssd1 vccd1 vccd1 _1806_/B sky130_fd_sc_hd__nor2_1
X_1734_ _1734_/A vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__clkbuf_2
X_1665_ _2114_/A _1795_/A _1665_/C _1665_/D vssd1 vssd1 vccd1 vccd1 _1666_/B sky130_fd_sc_hd__and4_1
X_1596_ _1593_/B _1595_/X _2498_/Q vssd1 vssd1 vccd1 vccd1 _1597_/C sky130_fd_sc_hd__a21oi_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2217_ _2221_/A vssd1 vssd1 vccd1 vccd1 _2217_/Y sky130_fd_sc_hd__inv_2
X_2079_ _2085_/A vssd1 vssd1 vccd1 vccd1 _2084_/A sky130_fd_sc_hd__buf_6
X_2148_ _2166_/A vssd1 vssd1 vccd1 vccd1 _2153_/A sky130_fd_sc_hd__buf_2
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1450_ _1450_/A vssd1 vssd1 vccd1 vccd1 _2528_/D sky130_fd_sc_hd__clkbuf_1
X_1381_ _1381_/A vssd1 vssd1 vccd1 vccd1 _2540_/D sky130_fd_sc_hd__inv_2
X_2002_ _2004_/A vssd1 vssd1 vccd1 vccd1 _2002_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2766_ _2766_/A _2068_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_2697_ _2697_/A _1985_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_1717_ _2473_/Q _1703_/X _1715_/X _1716_/X vssd1 vssd1 vccd1 vccd1 _2473_/D sky130_fd_sc_hd__a22o_1
X_1648_ _1645_/Y _1650_/B _1647_/X vssd1 vssd1 vccd1 vccd1 _2483_/D sky130_fd_sc_hd__a21oi_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1579_/A vssd1 vssd1 vccd1 vccd1 _2504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2551_ _2560_/CLK _2551_/D vssd1 vssd1 vccd1 vccd1 _2551_/Q sky130_fd_sc_hd__dfxtp_1
X_2482_ _2544_/CLK _2482_/D _2215_/Y vssd1 vssd1 vccd1 vccd1 _2482_/Q sky130_fd_sc_hd__dfrtp_1
X_1502_ _1513_/A vssd1 vssd1 vccd1 vccd1 _1503_/B sky130_fd_sc_hd__buf_2
X_1433_ _1474_/A _1433_/B vssd1 vssd1 vccd1 vccd1 _1457_/B sky130_fd_sc_hd__nor2_2
X_1295_ _2510_/Q _2509_/Q _2480_/Q _2479_/Q vssd1 vssd1 vccd1 vccd1 _1298_/B sky130_fd_sc_hd__or4_1
X_1364_ _2533_/Q vssd1 vssd1 vccd1 vccd1 _1430_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2654__82 vssd1 vssd1 vccd1 vccd1 _2654__82/HI _2762_/A sky130_fd_sc_hd__conb_1
X_2749_ _2749_/A _2092_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1982_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1982_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2534_ _2537_/CLK _2534_/D _2279_/Y vssd1 vssd1 vccd1 vccd1 _2534_/Q sky130_fd_sc_hd__dfrtp_1
X_2465_ _2559_/CLK _2465_/D _2194_/Y vssd1 vssd1 vccd1 vccd1 _2465_/Q sky130_fd_sc_hd__dfrtp_1
X_2396_ _2393_/A _2407_/D _2403_/A vssd1 vssd1 vccd1 vccd1 _2396_/Y sky130_fd_sc_hd__o21ai_1
X_1416_ _1416_/A vssd1 vssd1 vccd1 vccd1 _1658_/A sky130_fd_sc_hd__buf_2
X_1347_ _1671_/A _1403_/A _1413_/A _1419_/A vssd1 vssd1 vccd1 vccd1 _1384_/B sky130_fd_sc_hd__and4_1
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1278_ _1519_/A _1519_/B _1278_/C _1278_/D vssd1 vssd1 vccd1 vccd1 _1278_/X sky130_fd_sc_hd__or4_4
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ _2252_/A vssd1 vssd1 vccd1 vccd1 _2250_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2181_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2181_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2624__52 vssd1 vssd1 vccd1 vccd1 _2624__52/HI _2732_/A sky130_fd_sc_hd__conb_1
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1965_ _1967_/A vssd1 vssd1 vccd1 vccd1 _1965_/Y sky130_fd_sc_hd__inv_2
X_1896_ _1341_/X _1897_/C _1824_/X vssd1 vssd1 vccd1 vccd1 _1896_/X sky130_fd_sc_hd__a21o_1
X_2517_ _2526_/CLK _2517_/D _2258_/Y vssd1 vssd1 vccd1 vccd1 _2517_/Q sky130_fd_sc_hd__dfrtp_1
X_2448_ _2476_/CLK _2448_/D _2174_/Y vssd1 vssd1 vccd1 vccd1 _2448_/Q sky130_fd_sc_hd__dfrtp_1
X_2379_ _2378_/X _2376_/Y _2566_/Q vssd1 vssd1 vccd1 vccd1 _2380_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1750_ _1754_/A _1757_/A _2466_/Q vssd1 vssd1 vccd1 vccd1 _1751_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1681_ _2448_/Q _2447_/Q _2446_/Q _2445_/Q vssd1 vssd1 vccd1 vccd1 _1812_/A sky130_fd_sc_hd__and4_1
X_2678__106 vssd1 vssd1 vccd1 vccd1 _2678__106/HI _2786_/A sky130_fd_sc_hd__conb_1
X_2164_ _2165_/A vssd1 vssd1 vccd1 vccd1 _2164_/Y sky130_fd_sc_hd__inv_2
X_2302_ _2302_/A vssd1 vssd1 vccd1 vccd1 _2302_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2233_ _2233_/A vssd1 vssd1 vccd1 vccd1 _2233_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2095_ _2407_/C vssd1 vssd1 vccd1 vccd1 _2302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1879_ _1876_/X _1878_/Y _2435_/Q vssd1 vssd1 vccd1 vccd1 _1880_/A sky130_fd_sc_hd__mux2_1
X_1948_ _2416_/Q _1947_/Y _1943_/X vssd1 vssd1 vccd1 vccd1 _2416_/D sky130_fd_sc_hd__o21a_1
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1802_ _2449_/Q _1812_/A vssd1 vssd1 vccd1 vccd1 _1803_/B sky130_fd_sc_hd__nand2_1
X_1733_ _1732_/A _1703_/X _1715_/X _1732_/Y vssd1 vssd1 vccd1 vccd1 _2470_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2782_ _2782_/A _2087_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664_ _1848_/A vssd1 vssd1 vccd1 vccd1 _1795_/A sky130_fd_sc_hd__buf_2
X_1595_ _1595_/A vssd1 vssd1 vccd1 vccd1 _1595_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2147_ _2147_/A vssd1 vssd1 vccd1 vccd1 _2147_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2216_ _2228_/A vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__buf_2
X_2078_ _2078_/A vssd1 vssd1 vccd1 vccd1 _2078_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1380_ _1380_/A _1380_/B vssd1 vssd1 vccd1 vccd1 _1381_/A sky130_fd_sc_hd__or2_1
X_2001_ _2004_/A vssd1 vssd1 vccd1 vccd1 _2001_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1716_ _2473_/Q _1716_/B vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__xor2_1
X_2696_ _2696_/A _1984_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
X_2765_ _2765_/A _2066_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
XFILLER_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1647_ _1547_/X _1639_/C _1657_/A vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__a21o_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1577_/X _1574_/Y _1578_/S vssd1 vssd1 vccd1 vccd1 _1579_/A sky130_fd_sc_hd__mux2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2585__13 vssd1 vssd1 vccd1 vccd1 _2585__13/HI _2689_/A sky130_fd_sc_hd__conb_1
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _2574_/CLK _2550_/D vssd1 vssd1 vccd1 vccd1 _2550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2481_ _2544_/CLK _2481_/D _2214_/Y vssd1 vssd1 vccd1 vccd1 _2481_/Q sky130_fd_sc_hd__dfrtp_1
X_1501_ _1501_/A _1501_/B vssd1 vssd1 vccd1 vccd1 _1507_/A sky130_fd_sc_hd__nand2_1
X_1432_ _1432_/A vssd1 vssd1 vccd1 vccd1 _2533_/D sky130_fd_sc_hd__inv_2
X_1363_ _2534_/Q vssd1 vssd1 vccd1 vccd1 _1668_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1294_ _2508_/Q _2507_/Q _2506_/Q _2505_/Q vssd1 vssd1 vccd1 vccd1 _1298_/A sky130_fd_sc_hd__or4_1
X_2748_ _2748_/A _2047_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_2679_ _2679_/A _1963_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1981_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1986_/A sky130_fd_sc_hd__buf_6
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2533_ _2572_/CLK _2533_/D _2278_/Y vssd1 vssd1 vccd1 vccd1 _2533_/Q sky130_fd_sc_hd__dfrtp_1
X_2464_ _2464_/CLK _2464_/D _2193_/Y vssd1 vssd1 vccd1 vccd1 _2464_/Q sky130_fd_sc_hd__dfrtp_1
X_1415_ _1415_/A _1433_/B vssd1 vssd1 vccd1 vccd1 _1416_/A sky130_fd_sc_hd__or2_2
X_2395_ _2395_/A vssd1 vssd1 vccd1 vccd1 _2570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1346_ _2535_/Q vssd1 vssd1 vccd1 vccd1 _1419_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1277_ _1277_/A _1277_/B _1409_/A _1277_/D vssd1 vssd1 vccd1 vccd1 _1278_/D sky130_fd_sc_hd__or4_1
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2180_ _2184_/A vssd1 vssd1 vccd1 vccd1 _2180_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _1967_/A vssd1 vssd1 vccd1 vccd1 _1964_/Y sky130_fd_sc_hd__inv_2
X_1895_ _2430_/Q _1902_/A _1905_/A vssd1 vssd1 vccd1 vccd1 _1897_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2447_ _2476_/CLK _2447_/D _2171_/Y vssd1 vssd1 vccd1 vccd1 _2447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2516_ _2526_/CLK _2516_/D _2257_/Y vssd1 vssd1 vccd1 vccd1 _2516_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1329_ _2436_/Q _2430_/Q _2431_/Q _2437_/Q vssd1 vssd1 vccd1 vccd1 _1339_/A sky130_fd_sc_hd__or4bb_1
X_2378_ _2565_/Q _2378_/B vssd1 vssd1 vccd1 vccd1 _2378_/X sky130_fd_sc_hd__and2_1
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1680_ _1737_/B vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__clkbuf_2
X_2301_ _2301_/A _2301_/B _2301_/C vssd1 vssd1 vccd1 vccd1 _2301_/Y sky130_fd_sc_hd__nand3_1
X_2163_ _2165_/A vssd1 vssd1 vccd1 vccd1 _2163_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2232_ _2233_/A vssd1 vssd1 vccd1 vccd1 _2232_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2094_ input2/X _2094_/B vssd1 vssd1 vccd1 vccd1 _2407_/C sky130_fd_sc_hd__nor2_2
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1878_ _1878_/A _1878_/B vssd1 vssd1 vccd1 vccd1 _1878_/Y sky130_fd_sc_hd__nand2_1
X_1947_ _1947_/A _1947_/B vssd1 vssd1 vccd1 vccd1 _1947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1801_ _2450_/Q vssd1 vssd1 vccd1 vccd1 _1803_/A sky130_fd_sc_hd__inv_2
X_1732_ _1732_/A _1732_/B vssd1 vssd1 vccd1 vccd1 _1732_/Y sky130_fd_sc_hd__xnor2_1
X_1663_ _2114_/A _2727_/A _1743_/B vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__a21bo_1
X_2781_ _2781_/A _2086_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _2499_/Q _1597_/B _1590_/Y vssd1 vssd1 vccd1 vccd1 _2499_/D sky130_fd_sc_hd__o21a_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2146_ _2147_/A vssd1 vssd1 vccd1 vccd1 _2146_/Y sky130_fd_sc_hd__inv_2
X_2215_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2215_/Y sky130_fd_sc_hd__inv_2
X_2077_ _2078_/A vssd1 vssd1 vccd1 vccd1 _2077_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _2004_/A vssd1 vssd1 vccd1 vccd1 _2000_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2764_ _2764_/A _2065_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
X_1715_ _1715_/A vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__buf_2
X_1646_ _1654_/C _1646_/B vssd1 vssd1 vccd1 vccd1 _1650_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2695_ _2695_/A _1983_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _1589_/A _1577_/B _1577_/C vssd1 vssd1 vccd1 vccd1 _1577_/X sky130_fd_sc_hd__and3_1
X_2129_ _2290_/A vssd1 vssd1 vccd1 vccd1 _2134_/A sky130_fd_sc_hd__buf_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2544_/CLK _2480_/D _2213_/Y vssd1 vssd1 vccd1 vccd1 _2480_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1500_ _1493_/A _1493_/B _1497_/Y vssd1 vssd1 vccd1 vccd1 _2515_/D sky130_fd_sc_hd__o21a_1
X_1293_ _1278_/X _1289_/X _2290_/A vssd1 vssd1 vccd1 vccd1 _1293_/Y sky130_fd_sc_hd__o21ai_1
X_1431_ _1430_/Y _1430_/A _1431_/S vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__mux2_1
X_1362_ _1455_/A _1455_/B _1362_/C _1468_/C vssd1 vssd1 vccd1 vccd1 _1434_/A sky130_fd_sc_hd__and4_1
XFILLER_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2747_ _2747_/A _2046_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
X_1629_ _2484_/Q vssd1 vssd1 vccd1 vccd1 _1639_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2645__73 vssd1 vssd1 vccd1 vccd1 _2645__73/HI _2753_/A sky130_fd_sc_hd__conb_1
XFILLER_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1980_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1980_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2463_ _2560_/CLK _2463_/D _2192_/Y vssd1 vssd1 vccd1 vccd1 _2463_/Q sky130_fd_sc_hd__dfrtp_2
X_2532_ _2537_/CLK _2532_/D _2276_/Y vssd1 vssd1 vccd1 vccd1 _2532_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2394_ _2393_/Y _2391_/A _2570_/Q vssd1 vssd1 vccd1 vccd1 _2395_/A sky130_fd_sc_hd__mux2_1
X_1414_ _1519_/A _1409_/X _1414_/C _1414_/D vssd1 vssd1 vccd1 vccd1 _1433_/B sky130_fd_sc_hd__and4bb_1
X_1276_ _2520_/Q _1493_/A _1498_/S _2519_/Q vssd1 vssd1 vccd1 vccd1 _1277_/D sky130_fd_sc_hd__or4bb_1
X_1345_ _2536_/Q vssd1 vssd1 vccd1 vccd1 _1413_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2574_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1894_ _1906_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1905_/A sky130_fd_sc_hd__and2_1
X_1963_ _1967_/A vssd1 vssd1 vccd1 vccd1 _1963_/Y sky130_fd_sc_hd__inv_2
X_2446_ _2476_/CLK _2446_/D _2170_/Y vssd1 vssd1 vccd1 vccd1 _2446_/Q sky130_fd_sc_hd__dfrtp_1
X_2515_ _2526_/CLK _2515_/D _2256_/Y vssd1 vssd1 vccd1 vccd1 _2515_/Q sky130_fd_sc_hd__dfrtp_1
X_1328_ _1710_/A vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__clkbuf_2
X_2377_ _2565_/Q _2378_/B _2376_/Y vssd1 vssd1 vccd1 vccd1 _2565_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1259_ _1259_/A vssd1 vssd1 vccd1 vccd1 _1492_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2615__43 vssd1 vssd1 vccd1 vccd1 _2615__43/HI _2719_/A sky130_fd_sc_hd__conb_1
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2300_ _2295_/X _2297_/Y _2298_/X _2299_/X _2301_/A vssd1 vssd1 vccd1 vccd1 _2546_/D
+ sky130_fd_sc_hd__a32o_1
X_2231_ _2233_/A vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__inv_2
X_2093_ _2093_/A vssd1 vssd1 vccd1 vccd1 _2093_/Y sky130_fd_sc_hd__inv_2
X_2162_ _2165_/A vssd1 vssd1 vccd1 vccd1 _2162_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1877_ _2434_/Q _2433_/Q _1885_/B _1886_/A vssd1 vssd1 vccd1 vccd1 _1878_/B sky130_fd_sc_hd__a31o_1
X_1946_ _1946_/A vssd1 vssd1 vccd1 vccd1 _1947_/B sky130_fd_sc_hd__inv_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2429_ _2431_/CLK _2429_/D _2150_/Y vssd1 vssd1 vccd1 vccd1 _2429_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1800_ _1800_/A vssd1 vssd1 vccd1 vccd1 _1800_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1731_ _1731_/A vssd1 vssd1 vccd1 vccd1 _2471_/D sky130_fd_sc_hd__clkbuf_1
X_1662_ _1662_/A vssd1 vssd1 vccd1 vccd1 _1743_/B sky130_fd_sc_hd__clkbuf_2
X_2780_ _2780_/A _2084_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
XFILLER_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2214_/Y sky130_fd_sc_hd__inv_2
X_1593_ _2498_/Q _1593_/B _1593_/C vssd1 vssd1 vccd1 vccd1 _1597_/B sky130_fd_sc_hd__and3_1
X_2145_ _2147_/A vssd1 vssd1 vccd1 vccd1 _2145_/Y sky130_fd_sc_hd__inv_2
X_2076_ _2078_/A vssd1 vssd1 vccd1 vccd1 _2076_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1929_ _2421_/Q _1923_/Y _1928_/Y _1924_/X _2422_/Q vssd1 vssd1 vccd1 vccd1 _2422_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2491_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2763_ _2763_/A _2064_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_1714_ _1734_/A vssd1 vssd1 vccd1 vccd1 _1715_/A sky130_fd_sc_hd__clkbuf_2
X_1645_ _2483_/Q vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__inv_2
X_1576_ _1573_/Y _1574_/Y _1575_/X vssd1 vssd1 vccd1 vccd1 _2505_/D sky130_fd_sc_hd__o21a_1
X_2694_ _2694_/A _1982_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2128_ _2128_/A vssd1 vssd1 vccd1 vccd1 _2411_/D sky130_fd_sc_hd__clkbuf_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2060_/A vssd1 vssd1 vccd1 vccd1 _2059_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1430_ _1430_/A _1650_/A vssd1 vssd1 vccd1 vccd1 _1430_/Y sky130_fd_sc_hd__nand2_1
X_1292_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2290_/A sky130_fd_sc_hd__buf_2
X_1361_ _2522_/Q _1472_/A _2520_/Q _2519_/Q vssd1 vssd1 vccd1 vccd1 _1468_/C sky130_fd_sc_hd__and4_1
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2746_ _2746_/A _2045_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
X_1628_ _1637_/A _1628_/B _1628_/C vssd1 vssd1 vccd1 vccd1 _2488_/D sky130_fd_sc_hd__nor3_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1559_ _1559_/A vssd1 vssd1 vccd1 vccd1 _1589_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660__88 vssd1 vssd1 vccd1 vccd1 _2660__88/HI _2768_/A sky130_fd_sc_hd__conb_1
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2462_ _2560_/CLK _2462_/D _2190_/Y vssd1 vssd1 vccd1 vccd1 _2462_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2393_ _2393_/A _2393_/B vssd1 vssd1 vccd1 vccd1 _2393_/Y sky130_fd_sc_hd__nor2_1
X_2531_ _2537_/CLK _2531_/D _2275_/Y vssd1 vssd1 vccd1 vccd1 _2531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1413_ _1413_/A _1413_/B _2526_/Q _1457_/A vssd1 vssd1 vccd1 vccd1 _1414_/D sky130_fd_sc_hd__and4_1
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1275_ _2516_/Q vssd1 vssd1 vccd1 vccd1 _1498_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_1344_ _2537_/Q vssd1 vssd1 vccd1 vccd1 _1403_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2729_ _2729_/A _2023_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _2093_/A vssd1 vssd1 vccd1 vccd1 _1967_/A sky130_fd_sc_hd__buf_8
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1893_ _2429_/Q vssd1 vssd1 vccd1 vccd1 _1902_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2445_ _2476_/CLK _2445_/D _2169_/Y vssd1 vssd1 vccd1 vccd1 _2445_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2376_ _2403_/A _2376_/B vssd1 vssd1 vccd1 vccd1 _2376_/Y sky130_fd_sc_hd__nand2_1
X_2514_ _2566_/CLK _2514_/D _2255_/Y vssd1 vssd1 vccd1 vccd1 _2514_/Q sky130_fd_sc_hd__dfrtp_1
X_1327_ _1665_/C _1665_/D _1304_/Y vssd1 vssd1 vccd1 vccd1 _1710_/A sky130_fd_sc_hd__a21o_1
X_1258_ _2544_/Q _1387_/B vssd1 vssd1 vccd1 vccd1 _1259_/A sky130_fd_sc_hd__and2_1
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2630__58 vssd1 vssd1 vccd1 vccd1 _2630__58/HI _2738_/A sky130_fd_sc_hd__conb_1
XFILLER_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2230_ _2233_/A vssd1 vssd1 vccd1 vccd1 _2230_/Y sky130_fd_sc_hd__inv_2
X_2161_ _2165_/A vssd1 vssd1 vccd1 vccd1 _2161_/Y sky130_fd_sc_hd__inv_2
X_2092_ _2093_/A vssd1 vssd1 vccd1 vccd1 _2092_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1945_ _2417_/Q _1943_/X _1944_/Y _1307_/X vssd1 vssd1 vccd1 vccd1 _2417_/D sky130_fd_sc_hd__a22o_1
X_1876_ _2434_/Q _2433_/Q _1916_/A _1885_/B vssd1 vssd1 vccd1 vccd1 _1876_/X sky130_fd_sc_hd__and4_1
X_2428_ _2431_/CLK _2428_/D _2149_/Y vssd1 vssd1 vccd1 vccd1 _2428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2359_ _2374_/C vssd1 vssd1 vccd1 vccd1 _2382_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1730_ _1730_/A _1730_/B vssd1 vssd1 vccd1 vccd1 _1731_/A sky130_fd_sc_hd__and2_1
X_1661_ _1659_/A _1625_/A _1660_/X vssd1 vssd1 vccd1 vccd1 _2479_/D sky130_fd_sc_hd__a21oi_1
XFILLER_7_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1592_ _1592_/A vssd1 vssd1 vccd1 vccd1 _2500_/D sky130_fd_sc_hd__clkbuf_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _2147_/A vssd1 vssd1 vccd1 vccd1 _2144_/Y sky130_fd_sc_hd__inv_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2213_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2213_/Y sky130_fd_sc_hd__inv_2
X_2075_ _2078_/A vssd1 vssd1 vccd1 vccd1 _2075_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1859_ _2423_/Q vssd1 vssd1 vccd1 vccd1 _1925_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1928_ _1928_/A _1928_/B vssd1 vssd1 vccd1 vccd1 _1928_/Y sky130_fd_sc_hd__nor2_1
X_2600__28 vssd1 vssd1 vccd1 vccd1 _2600__28/HI _2704_/A sky130_fd_sc_hd__conb_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2666__94 vssd1 vssd1 vccd1 vccd1 _2666__94/HI _2774_/A sky130_fd_sc_hd__conb_1
X_1713_ _1742_/A vssd1 vssd1 vccd1 vccd1 _1734_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2762_ _2762_/A _2063_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_2693_ _2693_/A _1980_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_1644_ _1644_/A vssd1 vssd1 vccd1 vccd1 _2484_/D sky130_fd_sc_hd__clkbuf_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ _1578_/S _1547_/X _1577_/C _2505_/Q vssd1 vssd1 vccd1 vccd1 _1575_/X sky130_fd_sc_hd__a31o_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _2126_/Y _2121_/A _2411_/Q vssd1 vssd1 vccd1 vccd1 _2128_/A sky130_fd_sc_hd__mux2_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2058_ _2060_/A vssd1 vssd1 vccd1 vccd1 _2058_/Y sky130_fd_sc_hd__inv_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1360_ _2521_/Q vssd1 vssd1 vccd1 vccd1 _1472_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2591__19 vssd1 vssd1 vccd1 vccd1 _2591__19/HI _2695_/A sky130_fd_sc_hd__conb_1
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1291_ _2234_/A vssd1 vssd1 vccd1 vccd1 _2283_/A sky130_fd_sc_hd__buf_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2745_ _2745_/A _2044_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1627_ _1634_/A _1634_/B _2488_/Q vssd1 vssd1 vccd1 vccd1 _1628_/C sky130_fd_sc_hd__a21oi_1
X_1558_ _2508_/Q _1554_/X _1555_/Y _1625_/A vssd1 vssd1 vccd1 vccd1 _2508_/D sky130_fd_sc_hd__a22o_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _1402_/X _1484_/Y _1488_/X vssd1 vssd1 vccd1 vccd1 _2518_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2636__64 vssd1 vssd1 vccd1 vccd1 _2636__64/HI _2744_/A sky130_fd_sc_hd__conb_1
X_2530_ _2537_/CLK _2530_/D _2274_/Y vssd1 vssd1 vccd1 vccd1 _2530_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2461_ _2560_/CLK _2461_/D _2189_/Y vssd1 vssd1 vccd1 vccd1 _2461_/Q sky130_fd_sc_hd__dfrtp_1
X_2392_ _2392_/A vssd1 vssd1 vccd1 vccd1 _2569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1412_ _2535_/Q vssd1 vssd1 vccd1 vccd1 _1413_/B sky130_fd_sc_hd__inv_2
X_1343_ _2538_/Q vssd1 vssd1 vccd1 vccd1 _1671_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1274_ _2515_/Q vssd1 vssd1 vccd1 vccd1 _1493_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2728_ input2/X _2022_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ _2085_/A vssd1 vssd1 vccd1 vccd1 _2093_/A sky130_fd_sc_hd__buf_8
X_1892_ _1892_/A vssd1 vssd1 vccd1 vccd1 _2432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2513_ _2566_/CLK _2513_/D _2254_/Y vssd1 vssd1 vccd1 vccd1 _2513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2444_ _2559_/CLK _2444_/D _2168_/Y vssd1 vssd1 vccd1 vccd1 _2725_/A sky130_fd_sc_hd__dfrtp_2
X_1326_ _2113_/B _2113_/C _1662_/A vssd1 vssd1 vccd1 vccd1 _2094_/B sky130_fd_sc_hd__a21o_1
X_2375_ _2382_/A _2565_/Q _2372_/C _2393_/A vssd1 vssd1 vccd1 vccd1 _2376_/B sky130_fd_sc_hd__a31o_1
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1257_ _2543_/Q vssd1 vssd1 vccd1 vccd1 _1387_/B sky130_fd_sc_hd__inv_2
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2606__34 vssd1 vssd1 vccd1 vccd1 _2606__34/HI _2710_/A sky130_fd_sc_hd__conb_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2160_ _2166_/A vssd1 vssd1 vccd1 vccd1 _2165_/A sky130_fd_sc_hd__buf_2
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2091_ _2093_/A vssd1 vssd1 vccd1 vccd1 _2091_/Y sky130_fd_sc_hd__inv_2
X_1875_ _2432_/Q _1875_/B _1906_/B vssd1 vssd1 vccd1 vccd1 _1885_/B sky130_fd_sc_hd__and3_1
X_1944_ _2417_/Q _1944_/B vssd1 vssd1 vccd1 vccd1 _1944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2427_ _2431_/CLK _2427_/D _2147_/Y vssd1 vssd1 vccd1 vccd1 _2427_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2289_ _2290_/A vssd1 vssd1 vccd1 vccd1 _2289_/Y sky130_fd_sc_hd__inv_2
X_1309_ _2544_/Q vssd1 vssd1 vccd1 vccd1 _1387_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2358_ _2561_/Q _2358_/B _2358_/C vssd1 vssd1 vccd1 vccd1 _2374_/C sky130_fd_sc_hd__and3_1
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _1474_/X _1278_/X _1658_/Y _1659_/Y vssd1 vssd1 vccd1 vccd1 _1660_/X sky130_fd_sc_hd__o31a_1
X_1591_ _1589_/X _1590_/Y _1591_/S vssd1 vssd1 vccd1 vccd1 _1592_/A sky130_fd_sc_hd__mux2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _2147_/A vssd1 vssd1 vccd1 vccd1 _2143_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2212_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2212_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2074_ _2078_/A vssd1 vssd1 vccd1 vccd1 _2074_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2597__25 vssd1 vssd1 vccd1 vccd1 _2597__25/HI _2701_/A sky130_fd_sc_hd__conb_1
X_1927_ _2420_/Q _1933_/A vssd1 vssd1 vccd1 vccd1 _1928_/B sky130_fd_sc_hd__nand2_1
X_1858_ _1946_/A _1936_/C _1858_/C vssd1 vssd1 vccd1 vccd1 _1933_/A sky130_fd_sc_hd__and3_1
X_1789_ _1789_/A _1789_/B vssd1 vssd1 vccd1 vccd1 _1789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2692_ _2692_/A _1979_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1712_ _1886_/A _1743_/B _1712_/C vssd1 vssd1 vccd1 vccd1 _1742_/A sky130_fd_sc_hd__and3_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1643_ _1643_/A _1643_/B _1643_/C vssd1 vssd1 vccd1 vccd1 _1644_/A sky130_fd_sc_hd__and3_1
X_2761_ _2761_/A _2062_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _1474_/A _1577_/C _1639_/B vssd1 vssd1 vccd1 vccd1 _1574_/Y sky130_fd_sc_hd__o21ai_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _2386_/A _2126_/B vssd1 vssd1 vccd1 vccd1 _2126_/Y sky130_fd_sc_hd__nor2_1
X_2057_ _2060_/A vssd1 vssd1 vccd1 vccd1 _2057_/Y sky130_fd_sc_hd__inv_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2674__102 vssd1 vssd1 vccd1 vccd1 _2674__102/HI _2782_/A sky130_fd_sc_hd__conb_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1290_ input2/X vssd1 vssd1 vccd1 vccd1 _2234_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1626_ _2489_/Q _1628_/B _1625_/Y _1503_/B vssd1 vssd1 vccd1 vccd1 _2489_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2744_ _2744_/A _2042_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_1557_ _1633_/A vssd1 vssd1 vccd1 vccd1 _1625_/A sky130_fd_sc_hd__clkbuf_2
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _1455_/A _1487_/X _1457_/B _2518_/Q vssd1 vssd1 vccd1 vccd1 _1488_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2109_ _2557_/Q _2560_/Q _2109_/C _2109_/D vssd1 vssd1 vccd1 vccd1 _2358_/C sky130_fd_sc_hd__and4_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2651__79 vssd1 vssd1 vccd1 vccd1 _2651__79/HI _2759_/A sky130_fd_sc_hd__conb_1
X_2460_ _2560_/CLK _2460_/D _2188_/Y vssd1 vssd1 vccd1 vccd1 _2460_/Q sky130_fd_sc_hd__dfrtp_1
X_1342_ _1304_/Y _1312_/Y _2094_/B _1341_/X vssd1 vssd1 vccd1 vccd1 _2543_/D sky130_fd_sc_hd__a31o_1
X_2391_ _2391_/A _2391_/B vssd1 vssd1 vccd1 vccd1 _2392_/A sky130_fd_sc_hd__and2_1
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1411_ _2528_/Q _2523_/Q _1465_/A _1453_/A vssd1 vssd1 vccd1 vccd1 _1414_/C sky130_fd_sc_hd__and4bb_1
X_1273_ _2538_/Q _2537_/Q _2533_/Q _2534_/Q vssd1 vssd1 vccd1 vccd1 _1409_/A sky130_fd_sc_hd__or4b_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2727_ _2727_/A _2021_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
X_1609_ _1609_/A vssd1 vssd1 vccd1 vccd1 _2494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1960_ input1/X vssd1 vssd1 vccd1 vccd1 _2085_/A sky130_fd_sc_hd__buf_2
X_1891_ _1891_/A _1891_/B vssd1 vssd1 vccd1 vccd1 _1892_/A sky130_fd_sc_hd__and2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2443_ _2544_/CLK _2443_/D _2167_/Y vssd1 vssd1 vccd1 vccd1 _2443_/Q sky130_fd_sc_hd__dfrtp_1
X_2512_ _2568_/CLK _2512_/D _2252_/Y vssd1 vssd1 vccd1 vccd1 _2512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1325_ _1387_/A _1848_/A vssd1 vssd1 vccd1 vccd1 _1662_/A sky130_fd_sc_hd__or2_1
X_2374_ _2374_/A _2407_/C _2374_/C vssd1 vssd1 vccd1 vccd1 _2378_/B sky130_fd_sc_hd__and3_1
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2621__49 vssd1 vssd1 vccd1 vccd1 _2621__49/HI _2729_/A sky130_fd_sc_hd__conb_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2090_ _2090_/A vssd1 vssd1 vccd1 vccd1 _2090_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2572_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1874_ _2423_/Q _1874_/B _1908_/C vssd1 vssd1 vccd1 vccd1 _1906_/B sky130_fd_sc_hd__and3_1
X_1943_ _1307_/A _1944_/B _1903_/A vssd1 vssd1 vccd1 vccd1 _1943_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2426_ _2439_/CLK _2426_/D _2146_/Y vssd1 vssd1 vccd1 vccd1 _2426_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2357_ _2561_/Q _2357_/B vssd1 vssd1 vccd1 vccd1 _2357_/X sky130_fd_sc_hd__or2_1
X_1308_ _1501_/A _1293_/Y _1307_/X vssd1 vssd1 vccd1 vccd1 _2544_/D sky130_fd_sc_hd__a21o_1
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2288_ _2288_/A vssd1 vssd1 vccd1 vccd1 _2288_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _1589_/B _1595_/A _1569_/A vssd1 vssd1 vccd1 vccd1 _1590_/Y sky130_fd_sc_hd__a21oi_1
X_2073_ _2085_/A vssd1 vssd1 vccd1 vccd1 _2078_/A sky130_fd_sc_hd__buf_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _2166_/A vssd1 vssd1 vccd1 vccd1 _2147_/A sky130_fd_sc_hd__buf_2
X_2211_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2211_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1926_ _1925_/A _1924_/X _1925_/Y _1908_/C vssd1 vssd1 vccd1 vccd1 _2423_/D sky130_fd_sc_hd__a22o_1
X_1788_ _1788_/A _1788_/B vssd1 vssd1 vccd1 vccd1 _1789_/B sky130_fd_sc_hd__nor2_1
X_1857_ _1857_/A vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2409_ _2409_/A vssd1 vssd1 vccd1 vccd1 _2574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2691_ _2691_/A _1978_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
X_1711_ _2113_/A _1743_/C vssd1 vssd1 vccd1 vccd1 _1712_/C sky130_fd_sc_hd__and2_1
X_2760_ _2760_/A _2060_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
X_1642_ _1577_/B _1632_/A _1639_/A vssd1 vssd1 vccd1 vccd1 _1643_/C sky130_fd_sc_hd__a21o_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _2505_/Q _1578_/S _1555_/B vssd1 vssd1 vccd1 vccd1 _1573_/Y sky130_fd_sc_hd__a21oi_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2056_ _2060_/A vssd1 vssd1 vccd1 vccd1 _2056_/Y sky130_fd_sc_hd__inv_2
X_2125_ _2367_/A vssd1 vssd1 vccd1 vccd1 _2386_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2657__85 vssd1 vssd1 vccd1 vccd1 _2657__85/HI _2765_/A sky130_fd_sc_hd__conb_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1909_ _2426_/Q _2425_/Q _1916_/B vssd1 vssd1 vccd1 vccd1 _1909_/X sky130_fd_sc_hd__and3_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2743_ _2743_/A _2041_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1625_ _1625_/A _1625_/B vssd1 vssd1 vccd1 vccd1 _1625_/Y sky130_fd_sc_hd__nand2_1
X_1556_ _1612_/A vssd1 vssd1 vccd1 vccd1 _1633_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1670_/D _1498_/S _1493_/A vssd1 vssd1 vccd1 vccd1 _1487_/X sky130_fd_sc_hd__and3_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2108_ _2558_/Q _2559_/Q vssd1 vssd1 vccd1 vccd1 _2109_/D sky130_fd_sc_hd__and2_1
X_2039_ _2042_/A vssd1 vssd1 vccd1 vccd1 _2039_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2439_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1410_ _2527_/Q vssd1 vssd1 vccd1 vccd1 _1453_/A sky130_fd_sc_hd__clkbuf_1
X_1341_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1341_/X sky130_fd_sc_hd__buf_2
X_2390_ _2110_/B _2302_/A _2357_/B _2569_/Q vssd1 vssd1 vccd1 vccd1 _2391_/B sky130_fd_sc_hd__a31o_1
X_1272_ _2526_/Q _2521_/Q _2522_/Q _2525_/Q vssd1 vssd1 vccd1 vccd1 _1277_/B sky130_fd_sc_hd__or4bb_1
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2627__55 vssd1 vssd1 vccd1 vccd1 _2627__55/HI _2735_/A sky130_fd_sc_hd__conb_1
X_2726_ _2726_/A _2020_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
X_1608_ _1643_/A _1608_/B _1608_/C vssd1 vssd1 vccd1 vccd1 _1609_/A sky130_fd_sc_hd__and3_1
X_1539_ _1559_/A _1539_/B _1604_/B vssd1 vssd1 vccd1 vccd1 _1570_/B sky130_fd_sc_hd__and3_1
XFILLER_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1890_ _1885_/A _1875_/B _1906_/B _2432_/Q vssd1 vssd1 vccd1 vccd1 _1891_/B sky130_fd_sc_hd__a31o_1
X_2442_ _2544_/CLK _2442_/D _2165_/Y vssd1 vssd1 vccd1 vccd1 _2442_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2511_ _2568_/CLK _2511_/D _2251_/Y vssd1 vssd1 vccd1 vccd1 _2511_/Q sky130_fd_sc_hd__dfrtp_1
X_2373_ _2382_/A _2369_/Y _2372_/X vssd1 vssd1 vccd1 vccd1 _2564_/D sky130_fd_sc_hd__a21o_1
XFILLER_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1324_ _2543_/Q vssd1 vssd1 vccd1 vccd1 _1848_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _2709_/A _2000_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1942_ _2416_/Q _1946_/A vssd1 vssd1 vccd1 vccd1 _1944_/B sky130_fd_sc_hd__nand2_1
X_1873_ _1844_/X _2436_/Q _1871_/X _1872_/Y vssd1 vssd1 vccd1 vccd1 _2436_/D sky130_fd_sc_hd__a22o_1
X_2425_ _2439_/CLK _2425_/D _2145_/Y vssd1 vssd1 vccd1 vccd1 _2425_/Q sky130_fd_sc_hd__dfrtp_1
X_2356_ _2356_/A _2358_/C vssd1 vssd1 vccd1 vccd1 _2357_/B sky130_fd_sc_hd__and2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1307_ _1307_/A vssd1 vssd1 vccd1 vccd1 _1307_/X sky130_fd_sc_hd__buf_2
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2287_ _2288_/A vssd1 vssd1 vccd1 vccd1 _2287_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2228_/A vssd1 vssd1 vccd1 vccd1 _2215_/A sky130_fd_sc_hd__clkbuf_2
X_2072_ _2072_/A vssd1 vssd1 vccd1 vccd1 _2072_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2141_ _2234_/A vssd1 vssd1 vccd1 vccd1 _2166_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1925_ _1925_/A _1947_/A vssd1 vssd1 vccd1 vccd1 _1925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1787_ _1787_/A _1787_/B vssd1 vssd1 vccd1 vccd1 _1788_/B sky130_fd_sc_hd__and2_1
X_1856_ _2439_/Q vssd1 vssd1 vccd1 vccd1 _1856_/Y sky130_fd_sc_hd__inv_2
X_2339_ _2298_/X _2337_/Y _2338_/X _2320_/X _2555_/Q vssd1 vssd1 vccd1 vccd1 _2555_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2408_ _2407_/X _2405_/A _2574_/Q vssd1 vssd1 vccd1 vccd1 _2409_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2588__16 vssd1 vssd1 vccd1 vccd1 _2588__16/HI _2692_/A sky130_fd_sc_hd__conb_1
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1710_ _1710_/A _1710_/B vssd1 vssd1 vccd1 vccd1 _1886_/A sky130_fd_sc_hd__or2_1
X_1641_ _1638_/Y _1643_/B _1640_/X _1503_/B vssd1 vssd1 vccd1 vccd1 _2485_/D sky130_fd_sc_hd__o211a_1
X_1572_ _1637_/A _1572_/B _1571_/X vssd1 vssd1 vccd1 vccd1 _2506_/D sky130_fd_sc_hd__nor3b_1
X_2690_ _2690_/A _1977_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_6_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2124_ _2323_/B _2124_/B vssd1 vssd1 vccd1 vccd1 _2367_/A sky130_fd_sc_hd__nand2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2060_/A sky130_fd_sc_hd__buf_6
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1908_ _2424_/Q _1925_/A _1908_/C vssd1 vssd1 vccd1 vccd1 _1916_/B sky130_fd_sc_hd__and3_1
X_1839_ _1928_/A vssd1 vssd1 vccd1 vccd1 _1947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2742_ _2742_/A _2040_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_1624_ _2488_/Q _1654_/C _1634_/B vssd1 vssd1 vccd1 vccd1 _1628_/B sky130_fd_sc_hd__and3_1
X_1555_ _2508_/Q _1555_/B _1555_/C vssd1 vssd1 vccd1 vccd1 _1555_/Y sky130_fd_sc_hd__nor3_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2107_ _2554_/Q _2553_/Q _2556_/Q _2555_/Q vssd1 vssd1 vccd1 vccd1 _2109_/C sky130_fd_sc_hd__and4_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _1483_/Y _1484_/A _1451_/X _1485_/X vssd1 vssd1 vccd1 vccd1 _2519_/D sky130_fd_sc_hd__a31o_1
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2038_ _2042_/A vssd1 vssd1 vccd1 vccd1 _2038_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1340_ _1928_/A _1710_/B vssd1 vssd1 vccd1 vccd1 _1916_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1271_ _2536_/Q _2535_/Q _2531_/Q _2532_/Q vssd1 vssd1 vccd1 vccd1 _1277_/A sky130_fd_sc_hd__or4b_1
X_2725_ _2725_/A _2019_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_1538_ _1646_/B _1562_/C _1563_/B _1538_/D vssd1 vssd1 vccd1 vccd1 _1604_/B sky130_fd_sc_hd__and4_1
X_1607_ _1639_/B _1606_/X _2494_/Q vssd1 vssd1 vccd1 vccd1 _1608_/C sky130_fd_sc_hd__a21o_1
X_1469_ _1467_/Y _1467_/A _1476_/A vssd1 vssd1 vccd1 vccd1 _1470_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2510_ _2566_/CLK _2510_/D _2250_/Y vssd1 vssd1 vccd1 vccd1 _2510_/Q sky130_fd_sc_hd__dfrtp_1
X_2441_ _2544_/CLK _2441_/D _2164_/Y vssd1 vssd1 vccd1 vccd1 _2441_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1323_ _1323_/A _1323_/B _1323_/C _1323_/D vssd1 vssd1 vccd1 vccd1 _2113_/C sky130_fd_sc_hd__nor4_2
X_2372_ _2382_/A _2372_/B _2372_/C vssd1 vssd1 vccd1 vccd1 _2372_/X sky130_fd_sc_hd__and3b_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2708_ _2708_/A _1998_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_59_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1872_ _1947_/A _1872_/B vssd1 vssd1 vccd1 vccd1 _1872_/Y sky130_fd_sc_hd__nor2_1
X_1941_ _1307_/X _1939_/Y _1940_/X _2418_/Q _1903_/X vssd1 vssd1 vccd1 vccd1 _2418_/D
+ sky130_fd_sc_hd__a32o_1
X_2424_ _2439_/CLK _2424_/D _2144_/Y vssd1 vssd1 vccd1 vccd1 _2424_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1306_ _1847_/B vssd1 vssd1 vccd1 vccd1 _1307_/A sky130_fd_sc_hd__clkbuf_2
X_2355_ _2560_/Q _2352_/Y _2354_/X vssd1 vssd1 vccd1 vccd1 _2560_/D sky130_fd_sc_hd__a21o_1
X_2286_ _2288_/A vssd1 vssd1 vccd1 vccd1 _2286_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2140_/A vssd1 vssd1 vccd1 vccd1 _2140_/Y sky130_fd_sc_hd__inv_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2071_ _2072_/A vssd1 vssd1 vccd1 vccd1 _2071_/Y sky130_fd_sc_hd__inv_2
X_1924_ _1307_/A _1923_/Y _1903_/A vssd1 vssd1 vccd1 vccd1 _1924_/X sky130_fd_sc_hd__a21o_1
X_1855_ _1855_/A vssd1 vssd1 vccd1 vccd1 _2440_/D sky130_fd_sc_hd__clkbuf_1
X_1786_ _1785_/A _1761_/X _1708_/A _1785_/X vssd1 vssd1 vccd1 vccd1 _2457_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2338_ _2336_/A _2336_/B _2356_/A _2555_/Q vssd1 vssd1 vccd1 vccd1 _2338_/X sky130_fd_sc_hd__a31o_1
X_2407_ _2407_/A _2573_/Q _2407_/C _2407_/D vssd1 vssd1 vccd1 vccd1 _2407_/X sky130_fd_sc_hd__and4_1
X_2269_ _2270_/A vssd1 vssd1 vccd1 vccd1 _2269_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1640_ _1639_/A _1547_/X _1639_/C _1638_/A vssd1 vssd1 vccd1 vccd1 _1640_/X sky130_fd_sc_hd__a31o_1
X_1571_ _2505_/Q _1578_/S _1633_/A _1577_/C _2506_/Q vssd1 vssd1 vccd1 vccd1 _1571_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2123_ _2113_/B _2113_/C _1743_/B vssd1 vssd1 vccd1 vccd1 _2124_/B sky130_fd_sc_hd__a21oi_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2054_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2054_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1907_ _1307_/X _1905_/Y _1906_/X _1906_/A _1903_/X vssd1 vssd1 vccd1 vccd1 _2428_/D
+ sky130_fd_sc_hd__a32o_1
X_1838_ _2441_/Q _2440_/Q _1847_/C vssd1 vssd1 vccd1 vccd1 _1845_/B sky130_fd_sc_hd__and3_1
X_1769_ _2458_/Q vssd1 vssd1 vccd1 vccd1 _1773_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2648__76 vssd1 vssd1 vccd1 vccd1 _2648__76/HI _2756_/A sky130_fd_sc_hd__conb_1
XFILLER_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2662__90 vssd1 vssd1 vccd1 vccd1 _2662__90/HI _2770_/A sky130_fd_sc_hd__conb_1
X_2741_ _2741_/A _2039_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1623_ _1637_/A _1623_/B _1623_/C vssd1 vssd1 vccd1 vccd1 _2490_/D sky130_fd_sc_hd__nor3_1
X_1554_ _1501_/A _1555_/C _1547_/X vssd1 vssd1 vccd1 vccd1 _1554_/X sky130_fd_sc_hd__a21bo_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1465_/B _1484_/Y _1483_/A vssd1 vssd1 vccd1 vccd1 _1485_/X sky130_fd_sc_hd__o21a_1
.ends

