magic
tech sky130A
magscale 1 2
timestamp 1654523694
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 658 2128 38824 37584
<< metal2 >>
rect -10 39200 102 40000
rect 634 39200 746 40000
rect 1278 39200 1390 40000
rect 1922 39200 2034 40000
rect 2566 39200 2678 40000
rect 3854 39200 3966 40000
rect 4498 39200 4610 40000
rect 5142 39200 5254 40000
rect 5786 39200 5898 40000
rect 6430 39200 6542 40000
rect 7074 39200 7186 40000
rect 7718 39200 7830 40000
rect 9006 39200 9118 40000
rect 9650 39200 9762 40000
rect 10294 39200 10406 40000
rect 10938 39200 11050 40000
rect 11582 39200 11694 40000
rect 12226 39200 12338 40000
rect 12870 39200 12982 40000
rect 14158 39200 14270 40000
rect 14802 39200 14914 40000
rect 15446 39200 15558 40000
rect 16090 39200 16202 40000
rect 16734 39200 16846 40000
rect 17378 39200 17490 40000
rect 18022 39200 18134 40000
rect 19310 39200 19422 40000
rect 19954 39200 20066 40000
rect 20598 39200 20710 40000
rect 21242 39200 21354 40000
rect 21886 39200 21998 40000
rect 22530 39200 22642 40000
rect 23174 39200 23286 40000
rect 24462 39200 24574 40000
rect 25106 39200 25218 40000
rect 25750 39200 25862 40000
rect 26394 39200 26506 40000
rect 27038 39200 27150 40000
rect 27682 39200 27794 40000
rect 28326 39200 28438 40000
rect 29614 39200 29726 40000
rect 30258 39200 30370 40000
rect 30902 39200 31014 40000
rect 31546 39200 31658 40000
rect 32190 39200 32302 40000
rect 32834 39200 32946 40000
rect 33478 39200 33590 40000
rect 34766 39200 34878 40000
rect 35410 39200 35522 40000
rect 36054 39200 36166 40000
rect 36698 39200 36810 40000
rect 37342 39200 37454 40000
rect 37986 39200 38098 40000
rect 38630 39200 38742 40000
rect 39274 39200 39386 40000
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
<< obsm2 >>
rect 802 39144 1222 39200
rect 1446 39144 1866 39200
rect 2090 39144 2510 39200
rect 2734 39144 3798 39200
rect 4022 39144 4442 39200
rect 4666 39144 5086 39200
rect 5310 39144 5730 39200
rect 5954 39144 6374 39200
rect 6598 39144 7018 39200
rect 7242 39144 7662 39200
rect 7886 39144 8950 39200
rect 9174 39144 9594 39200
rect 9818 39144 10238 39200
rect 10462 39144 10882 39200
rect 11106 39144 11526 39200
rect 11750 39144 12170 39200
rect 12394 39144 12814 39200
rect 13038 39144 14102 39200
rect 14326 39144 14746 39200
rect 14970 39144 15390 39200
rect 15614 39144 16034 39200
rect 16258 39144 16678 39200
rect 16902 39144 17322 39200
rect 17546 39144 17966 39200
rect 18190 39144 19254 39200
rect 19478 39144 19898 39200
rect 20122 39144 20542 39200
rect 20766 39144 21186 39200
rect 21410 39144 21830 39200
rect 22054 39144 22474 39200
rect 22698 39144 23118 39200
rect 23342 39144 24406 39200
rect 24630 39144 25050 39200
rect 25274 39144 25694 39200
rect 25918 39144 26338 39200
rect 26562 39144 26982 39200
rect 27206 39144 27626 39200
rect 27850 39144 28270 39200
rect 28494 39144 29558 39200
rect 29782 39144 30202 39200
rect 30426 39144 30846 39200
rect 31070 39144 31490 39200
rect 31714 39144 32134 39200
rect 32358 39144 32778 39200
rect 33002 39144 33422 39200
rect 33646 39144 34710 39200
rect 34934 39144 35354 39200
rect 35578 39144 35998 39200
rect 36222 39144 36642 39200
rect 36866 39144 37286 39200
rect 37510 39144 37930 39200
rect 38154 39144 38574 39200
rect 664 856 38714 39144
rect 802 31 1222 856
rect 1446 31 1866 856
rect 2090 31 2510 856
rect 2734 31 3154 856
rect 3378 31 3798 856
rect 4022 31 4442 856
rect 4666 31 5730 856
rect 5954 31 6374 856
rect 6598 31 7018 856
rect 7242 31 7662 856
rect 7886 31 8306 856
rect 8530 31 8950 856
rect 9174 31 9594 856
rect 9818 31 10882 856
rect 11106 31 11526 856
rect 11750 31 12170 856
rect 12394 31 12814 856
rect 13038 31 13458 856
rect 13682 31 14102 856
rect 14326 31 14746 856
rect 14970 31 16034 856
rect 16258 31 16678 856
rect 16902 31 17322 856
rect 17546 31 17966 856
rect 18190 31 18610 856
rect 18834 31 19254 856
rect 19478 31 19898 856
rect 20122 31 21186 856
rect 21410 31 21830 856
rect 22054 31 22474 856
rect 22698 31 23118 856
rect 23342 31 23762 856
rect 23986 31 24406 856
rect 24630 31 25050 856
rect 25274 31 26338 856
rect 26562 31 26982 856
rect 27206 31 27626 856
rect 27850 31 28270 856
rect 28494 31 28914 856
rect 29138 31 29558 856
rect 29782 31 30202 856
rect 30426 31 31490 856
rect 31714 31 32134 856
rect 32358 31 32778 856
rect 33002 31 33422 856
rect 33646 31 34066 856
rect 34290 31 34710 856
rect 34934 31 35354 856
rect 35578 31 36642 856
rect 36866 31 37286 856
rect 37510 31 37930 856
rect 38154 31 38574 856
<< metal3 >>
rect 0 39388 800 39628
rect 0 38708 800 38948
rect 39200 38708 40000 38948
rect 39200 38028 40000 38268
rect 0 37348 800 37588
rect 39200 37348 40000 37588
rect 0 36668 800 36908
rect 39200 36668 40000 36908
rect 0 35988 800 36228
rect 39200 35988 40000 36228
rect 0 35308 800 35548
rect 39200 35308 40000 35548
rect 0 34628 800 34868
rect 39200 34628 40000 34868
rect 0 33948 800 34188
rect 0 33268 800 33508
rect 39200 33268 40000 33508
rect 39200 32588 40000 32828
rect 0 31908 800 32148
rect 39200 31908 40000 32148
rect 0 31228 800 31468
rect 39200 31228 40000 31468
rect 0 30548 800 30788
rect 39200 30548 40000 30788
rect 0 29868 800 30108
rect 39200 29868 40000 30108
rect 0 29188 800 29428
rect 39200 29188 40000 29428
rect 0 28508 800 28748
rect 0 27828 800 28068
rect 39200 27828 40000 28068
rect 39200 27148 40000 27388
rect 0 26468 800 26708
rect 39200 26468 40000 26708
rect 0 25788 800 26028
rect 39200 25788 40000 26028
rect 0 25108 800 25348
rect 39200 25108 40000 25348
rect 0 24428 800 24668
rect 39200 24428 40000 24668
rect 0 23748 800 23988
rect 39200 23748 40000 23988
rect 0 23068 800 23308
rect 0 22388 800 22628
rect 39200 22388 40000 22628
rect 39200 21708 40000 21948
rect 0 21028 800 21268
rect 39200 21028 40000 21268
rect 0 20348 800 20588
rect 39200 20348 40000 20588
rect 0 19668 800 19908
rect 39200 19668 40000 19908
rect 0 18988 800 19228
rect 39200 18988 40000 19228
rect 0 18308 800 18548
rect 39200 18308 40000 18548
rect 0 17628 800 17868
rect 0 16948 800 17188
rect 39200 16948 40000 17188
rect 39200 16268 40000 16508
rect 0 15588 800 15828
rect 39200 15588 40000 15828
rect 0 14908 800 15148
rect 39200 14908 40000 15148
rect 0 14228 800 14468
rect 39200 14228 40000 14468
rect 0 13548 800 13788
rect 39200 13548 40000 13788
rect 0 12868 800 13108
rect 39200 12868 40000 13108
rect 0 12188 800 12428
rect 0 11508 800 11748
rect 39200 11508 40000 11748
rect 39200 10828 40000 11068
rect 0 10148 800 10388
rect 39200 10148 40000 10388
rect 0 9468 800 9708
rect 39200 9468 40000 9708
rect 0 8788 800 9028
rect 39200 8788 40000 9028
rect 0 8108 800 8348
rect 39200 8108 40000 8348
rect 0 7428 800 7668
rect 39200 7428 40000 7668
rect 0 6748 800 6988
rect 0 6068 800 6308
rect 39200 6068 40000 6308
rect 39200 5388 40000 5628
rect 0 4708 800 4948
rect 39200 4708 40000 4948
rect 0 4028 800 4268
rect 39200 4028 40000 4268
rect 0 3348 800 3588
rect 39200 3348 40000 3588
rect 0 2668 800 2908
rect 39200 2668 40000 2908
rect 0 1988 800 2228
rect 39200 1988 40000 2228
rect 0 1308 800 1548
rect 0 628 800 868
rect 39200 628 40000 868
rect 39200 -52 40000 188
<< obsm3 >>
rect 880 38628 39120 38861
rect 800 38348 39200 38628
rect 800 37948 39120 38348
rect 800 37668 39200 37948
rect 880 37268 39120 37668
rect 800 36988 39200 37268
rect 880 36588 39120 36988
rect 800 36308 39200 36588
rect 880 35908 39120 36308
rect 800 35628 39200 35908
rect 880 35228 39120 35628
rect 800 34948 39200 35228
rect 880 34548 39120 34948
rect 800 34268 39200 34548
rect 880 33868 39200 34268
rect 800 33588 39200 33868
rect 880 33188 39120 33588
rect 800 32908 39200 33188
rect 800 32508 39120 32908
rect 800 32228 39200 32508
rect 880 31828 39120 32228
rect 800 31548 39200 31828
rect 880 31148 39120 31548
rect 800 30868 39200 31148
rect 880 30468 39120 30868
rect 800 30188 39200 30468
rect 880 29788 39120 30188
rect 800 29508 39200 29788
rect 880 29108 39120 29508
rect 800 28828 39200 29108
rect 880 28428 39200 28828
rect 800 28148 39200 28428
rect 880 27748 39120 28148
rect 800 27468 39200 27748
rect 800 27068 39120 27468
rect 800 26788 39200 27068
rect 880 26388 39120 26788
rect 800 26108 39200 26388
rect 880 25708 39120 26108
rect 800 25428 39200 25708
rect 880 25028 39120 25428
rect 800 24748 39200 25028
rect 880 24348 39120 24748
rect 800 24068 39200 24348
rect 880 23668 39120 24068
rect 800 23388 39200 23668
rect 880 22988 39200 23388
rect 800 22708 39200 22988
rect 880 22308 39120 22708
rect 800 22028 39200 22308
rect 800 21628 39120 22028
rect 800 21348 39200 21628
rect 880 20948 39120 21348
rect 800 20668 39200 20948
rect 880 20268 39120 20668
rect 800 19988 39200 20268
rect 880 19588 39120 19988
rect 800 19308 39200 19588
rect 880 18908 39120 19308
rect 800 18628 39200 18908
rect 880 18228 39120 18628
rect 800 17948 39200 18228
rect 880 17548 39200 17948
rect 800 17268 39200 17548
rect 880 16868 39120 17268
rect 800 16588 39200 16868
rect 800 16188 39120 16588
rect 800 15908 39200 16188
rect 880 15508 39120 15908
rect 800 15228 39200 15508
rect 880 14828 39120 15228
rect 800 14548 39200 14828
rect 880 14148 39120 14548
rect 800 13868 39200 14148
rect 880 13468 39120 13868
rect 800 13188 39200 13468
rect 880 12788 39120 13188
rect 800 12508 39200 12788
rect 880 12108 39200 12508
rect 800 11828 39200 12108
rect 880 11428 39120 11828
rect 800 11148 39200 11428
rect 800 10748 39120 11148
rect 800 10468 39200 10748
rect 880 10068 39120 10468
rect 800 9788 39200 10068
rect 880 9388 39120 9788
rect 800 9108 39200 9388
rect 880 8708 39120 9108
rect 800 8428 39200 8708
rect 880 8028 39120 8428
rect 800 7748 39200 8028
rect 880 7348 39120 7748
rect 800 7068 39200 7348
rect 880 6668 39200 7068
rect 800 6388 39200 6668
rect 880 5988 39120 6388
rect 800 5708 39200 5988
rect 800 5308 39120 5708
rect 800 5028 39200 5308
rect 880 4628 39120 5028
rect 800 4348 39200 4628
rect 880 3948 39120 4348
rect 800 3668 39200 3948
rect 880 3268 39120 3668
rect 800 2988 39200 3268
rect 880 2588 39120 2988
rect 800 2308 39200 2588
rect 880 1908 39120 2308
rect 800 1628 39200 1908
rect 880 1228 39200 1628
rect 800 948 39200 1228
rect 880 548 39120 948
rect 800 268 39200 548
rect 800 35 39120 268
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 7235 3843 19488 36821
rect 19968 3843 34848 36821
rect 35328 3843 35453 36821
<< labels >>
rlabel metal3 s 0 36668 800 36908 6 active
port 1 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 21886 39200 21998 40000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s -10 39200 102 40000 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 39200 33268 40000 33508 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 14802 39200 14914 40000 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 39200 35308 40000 35548 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 39200 3348 40000 3588 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 7718 39200 7830 40000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 9650 39200 9762 40000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 39200 12868 40000 13108 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 7074 39200 7186 40000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 5142 39200 5254 40000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 39200 8788 40000 9028 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 39274 39200 39386 40000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 39200 15588 40000 15828 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 30258 39200 30370 40000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 34766 39200 34878 40000 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 39200 25108 40000 25348 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 35410 39200 35522 40000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 22530 39200 22642 40000 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 39200 24428 40000 24668 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 39200 38028 40000 38268 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 39200 26468 40000 26708 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 6430 39200 6542 40000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal3 s 39200 22388 40000 22628 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal3 s 39200 11508 40000 11748 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal3 s 39200 10828 40000 11068 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal2 s 10938 39200 11050 40000 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal3 s 39200 1988 40000 2228 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 28326 39200 28438 40000 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal2 s 11582 39200 11694 40000 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal2 s 31546 0 31658 800 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 39200 16948 40000 17188 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 1278 39200 1390 40000 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal2 s 19954 39200 20066 40000 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal2 s 20598 39200 20710 40000 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal2 s 37986 0 38098 800 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 39200 31228 40000 31468 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal2 s 23174 39200 23286 40000 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal3 s 39200 25788 40000 26028 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal2 s 32834 39200 32946 40000 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal2 s 1922 39200 2034 40000 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 32834 0 32946 800 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal2 s 9006 39200 9118 40000 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 17628 800 17868 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal3 s 0 8788 800 9028 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 0 14228 800 14468 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 39200 -52 40000 188 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 0 25788 800 26028 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal3 s 39200 14228 40000 14468 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal2 s 10294 39200 10406 40000 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal2 s 8362 0 8474 800 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal3 s 39200 37348 40000 37588 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 39200 21708 40000 21948 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal3 s 0 6068 800 6308 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal3 s 39200 31908 40000 32148 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 0 33268 800 33508 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal3 s 39200 21028 40000 21268 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 36698 39200 36810 40000 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal2 s 37342 0 37454 800 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal2 s 26394 39200 26506 40000 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal2 s 32190 39200 32302 40000 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal3 s 39200 18308 40000 18548 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal2 s 21886 0 21998 800 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal2 s 29614 39200 29726 40000 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal2 s 30902 39200 31014 40000 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 13514 0 13626 800 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal3 s 39200 628 40000 868 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal2 s 5786 0 5898 800 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal3 s 0 11508 800 11748 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal3 s 0 37348 800 37588 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal3 s 39200 5388 40000 5628 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal3 s 39200 32588 40000 32828 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal3 s 39200 30548 40000 30788 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal2 s 12226 39200 12338 40000 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal3 s 39200 35988 40000 36228 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal3 s 0 34628 800 34868 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal3 s 39200 23748 40000 23988 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 18022 39200 18134 40000 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal2 s 37986 39200 38098 40000 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 0 15588 800 15828 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 0 12188 800 12428 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal3 s 39200 6068 40000 6308 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 39200 4708 40000 4948 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 12870 39200 12982 40000 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 25106 39200 25218 40000 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 19310 39200 19422 40000 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 14158 39200 14270 40000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 38630 39200 38742 40000 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 39200 7428 40000 7668 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 39200 2668 40000 2908 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 634 39200 746 40000 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 33478 39200 33590 40000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 39200 19668 40000 19908 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 15446 39200 15558 40000 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 16090 39200 16202 40000 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_data_out[0]
port 148 nsew signal bidirectional
rlabel metal3 s 39200 9468 40000 9708 6 la1_data_out[10]
port 149 nsew signal bidirectional
rlabel metal2 s 18022 0 18134 800 6 la1_data_out[11]
port 150 nsew signal bidirectional
rlabel metal3 s 39200 36668 40000 36908 6 la1_data_out[12]
port 151 nsew signal bidirectional
rlabel metal2 s 3854 39200 3966 40000 6 la1_data_out[13]
port 152 nsew signal bidirectional
rlabel metal2 s 21242 39200 21354 40000 6 la1_data_out[14]
port 153 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 154 nsew signal bidirectional
rlabel metal3 s 39200 13548 40000 13788 6 la1_data_out[16]
port 155 nsew signal bidirectional
rlabel metal3 s 39200 29188 40000 29428 6 la1_data_out[17]
port 156 nsew signal bidirectional
rlabel metal2 s 4498 39200 4610 40000 6 la1_data_out[18]
port 157 nsew signal bidirectional
rlabel metal3 s 39200 20348 40000 20588 6 la1_data_out[19]
port 158 nsew signal bidirectional
rlabel metal3 s 0 35988 800 36228 6 la1_data_out[1]
port 159 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 la1_data_out[20]
port 160 nsew signal bidirectional
rlabel metal3 s 39200 34628 40000 34868 6 la1_data_out[21]
port 161 nsew signal bidirectional
rlabel metal2 s 24462 39200 24574 40000 6 la1_data_out[22]
port 162 nsew signal bidirectional
rlabel metal2 s 9650 0 9762 800 6 la1_data_out[23]
port 163 nsew signal bidirectional
rlabel metal3 s 39200 14908 40000 15148 6 la1_data_out[24]
port 164 nsew signal bidirectional
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 165 nsew signal bidirectional
rlabel metal3 s 39200 4028 40000 4268 6 la1_data_out[26]
port 166 nsew signal bidirectional
rlabel metal3 s 0 38708 800 38948 6 la1_data_out[27]
port 167 nsew signal bidirectional
rlabel metal2 s 35410 0 35522 800 6 la1_data_out[28]
port 168 nsew signal bidirectional
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 169 nsew signal bidirectional
rlabel metal2 s 16734 0 16846 800 6 la1_data_out[2]
port 170 nsew signal bidirectional
rlabel metal3 s 39200 10148 40000 10388 6 la1_data_out[30]
port 171 nsew signal bidirectional
rlabel metal3 s 39200 38708 40000 38948 6 la1_data_out[31]
port 172 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[3]
port 173 nsew signal bidirectional
rlabel metal2 s 36698 0 36810 800 6 la1_data_out[4]
port 174 nsew signal bidirectional
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 175 nsew signal bidirectional
rlabel metal3 s 39200 16268 40000 16508 6 la1_data_out[6]
port 176 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 177 nsew signal bidirectional
rlabel metal3 s 39200 29868 40000 30108 6 la1_data_out[8]
port 178 nsew signal bidirectional
rlabel metal2 s 37342 39200 37454 40000 6 la1_data_out[9]
port 179 nsew signal bidirectional
rlabel metal2 s 39274 0 39386 800 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 36054 39200 36166 40000 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 2566 39200 2678 40000 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 17378 39200 17490 40000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 25750 39200 25862 40000 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 16734 39200 16846 40000 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 31546 39200 31658 40000 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 39200 8108 40000 8348 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 39200 27828 40000 28068 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 6748 800 6988 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 39200 27148 40000 27388 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 22530 0 22642 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 27682 39200 27794 40000 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 27038 39200 27150 40000 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 5786 39200 5898 40000 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 213 nsew ground input
rlabel metal3 s 39200 18988 40000 19228 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4032352
string GDS_FILE /openlane/designs/wrapped_cpr/runs/RUN_2022.06.06_13.53.06/results/finishing/wrapped_cpr.magic.gds
string GDS_START 532674
<< end >>

